`ifndef WYCHERPROOF_SECP384R1_SHA3384_SV
`define WYCHERPROOF_SECP384R1_SHA3384_SV
typedef struct packed {
  int           tc_id;
  logic         valid;  // 1: expected pass; 0: expected fail (zero/oversized)
  logic [383:0]  hash;
  logic [383:0] x;
  logic [383:0] y;
  logic [383:0] r;
  logic [383:0] s;
} ecdsa_vector_secp384r1_sha3384;

localparam int TEST_VECTORS_SECP384R1_SHA3384_NUM = 286;

ecdsa_vector_secp384r1_sha3384 test_vectors_secp384r1_sha3384 [] = '{
  '{1, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'hc0bb0ee1bffc6c7b74609ec20c460ec47f4d068f33d601870778e5e474860d77834d744db219e6abae9c32912907efd2},
  '{2, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{92, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c0000, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=50 s_len=48
  '{93, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'hf11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a10000},  // OUT_OF_RANGE r_len=48 s_len=50
  '{97, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c0500, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=50 s_len=48
  '{98, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'hf11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a10500},  // OUT_OF_RANGE r_len=48 s_len=50
  '{113, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // r=0
  '{114, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{117, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h36a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{118, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3d44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{119, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db4cc, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{120, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd3921},
  '{121, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0034a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db4, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{122, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h00a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{123, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h003f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39},
  '{124, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h0044f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{125, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=49 s_len=48
  '{126, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=48 s_len=49
  '{129, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // r=0
  '{130, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{131, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726b4f0fdd1ba4eeb869ab3182345a88754178a3e92aa12ddbf, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=49 s_len=48
  '{132, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019727262a62cdd1e08fc7ea7efcbeb447385e3db20bbd10888ad9, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=49 s_len=48
  '{133, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcb5bd125927577e395cc960276249d63649e6fb379fe68d912724fb039e84258bd66f58f03082026d561dad822b24bb4, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{134, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcb5bd125927577e395cc960276249d63649e6fb379fe68d8d9d59d322e1f7038158103414bb8c7a1c24df442ef777527, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{135, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcb5bd125927577e395cc960276249d63649e6fb379fe68d94b0f022e45b11479654ce7dcba5778abe875c16d55ed2241, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=49 s_len=48
  '{136, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=49 s_len=48
  '{137, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcb5bd125927577e395cc960276249d63649e6fb379fe68d912724fb039e84258bd66f58f03082026d561dad822b24bb4, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},
  '{138, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78874db51f73e84e472ce6a716df47684a2b3c004470826314},  // OUT_OF_RANGE r_len=48 s_len=49
  '{139, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78f8871a1b8b79f2887cb28bb24de619545163cd6ed6f8102e},  // OUT_OF_RANGE r_len=48 s_len=49
  '{140, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'hc0bb0ee1bffc6c7b74609ec20c460ec47f4d068f33d6018740159862804edf982b33669b69693f30c1b019265c42c65f},
  '{141, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'hc0bb0ee1bffc6c7b74609ec20c460ec47f4d068f33d6018778b24ae08c17b1b8d31958e920b897b5d4c3ffbb8f7d9cec},  // OUT_OF_RANGE r_len=48 s_len=49
  '{142, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'h3f44f11e400393848b9f613df3b9f13b80b2f970cc29fe78bfea679d7fb12067d4cc99649696c0cf3e4fe6d9a3bd39a1},  // OUT_OF_RANGE r_len=48 s_len=49
  '{143, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h34a42eda6d8a881c6a3369fd89db629c9b61904c86019726ed8db04fc617bda742990a70fcf7dfd92a9e2527dd4db44c, 384'hc0bb0ee1bffc6c7b74609ec20c460ec47f4d068f33d6018740159862804edf982b33669b69693f30c1b019265c42c65f},
  '{144, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // r=0, s=0
  '{145, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},  // r=0
  '{146, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},  // r=0
  '{147, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // r=0
  '{148, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // r=0
  '{149, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // r=0
  '{150, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // r=0
  '{151, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // r=0
  '{154, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{155, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{156, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{157, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{158, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{159, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{160, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{161, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{164, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{165, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{166, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{167, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{168, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{169, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{170, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{171, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{174, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{175, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{176, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{177, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{178, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{179, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{180, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{181, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{184, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{185, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{186, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{187, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{188, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{189, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{190, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{191, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{194, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{195, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{196, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{197, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{198, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{199, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{200, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{201, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{204, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{205, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{206, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{207, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{208, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{209, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{210, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{211, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{214, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{215, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{216, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{217, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{218, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{219, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{220, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{221, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{230, 1'b1, 384'hffcdf27e6dbfcd0798cb013f1240f6f1fd845a3d89ec16d3aad7ae298bfb1b13f7acdec4306f49346826cd80ac3adb76, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hac042e13ab83394692019170707bc21dd3d7b8d233d11b651757085bdd5767eabbb85322984f14437335de0cdf565684, 384'hc1045ed26ae9e8aabf5307db317f60e8c2842f67df81da26633d831ae5e061a5ef850d7d49f085d566d92cfd9f152d46},
  '{231, 1'b1, 384'h00000000d8f34863f5150caabbcdd0b014cb8f5e6c6215f81616752f6fdff77afb635307cb129730b5bcd1fe5f313564, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0c0b82be4c36d506063fc963133c14d5014d65c9eb796ee8a8387120119ccc16b57302b6ccb19a846b7762375b3c9718, 384'h285919259f684f56f89cbaa789ef13e185fd24d09dcd46ce794aedc4e5b4a3820535213abb7c4e605b02200fbeb3227c},
  '{232, 1'b1, 384'h9100000000d676979ba28b302bda3c58435097e95cf9385cff9de0096fd143fc32707bab8bc02c8ab981c0f7941c562a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7da99d7e8bb505cc5f12706d5eb7669336a61a726a5b376ff96d678a621f38681bc78592cd06717cb87753daf0d39b77, 384'hca91cdb78f21950877b69db1418a3e9b5799b3464f1fa223c7ac8d6fa9f647f2a08109935ad67477c96bbf1a2a127a1d},
  '{233, 1'b1, 384'ha4fa000000004b0fa23b91acb4ac09179f5a213e89d1f0b81972d8e88762c9b4319197336b136ab82a1d8edaa79fa1cd, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h204d322af7178ac20b39a42723fb1f8329b105993e09dbdcabf3e0eaa0a08d54719e06ba704691295a56be7765b5fd74, 384'h3b526de3e47e69518d4fbc0833a5785074c3f4eef27b9f0fc48481514931e43235b81e51d2b577b1739964ef25d8faad},
  '{234, 1'b1, 384'h6b142300000000b5b417c1787ce455d838edb8e8b55870b2c71ba7d0ab4fcd3c37e740f4a19755b26f5f92a04a90efd4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9d4adb54f52349cc73322ffc946bf44a1a1bb954bd4b58f912be068ce05272a12479bbb0f778a9faf8f9f2e9324bd5e9, 384'h1eee2f98406c30728da3b2b533c387108cc67fc24abdb6bdab686f207f0a75cc9c3b4d4ea9427d881c47d419ed7a1b95},
  '{235, 1'b1, 384'hfa5c4faa00000000aed513501d57b72424151f517517883e6a63f366bff660bdef8b655e5c4d45c77af93ef0f98bc3d8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hae50b1aaad54efbe007f1da7d50ec00cf1100f904fd8f4940ef48f364031dc1284ab984e018105e6d368bb5a47c25022, 384'ha803fb0156a10e42d4294a764a1da9c3e0c8320bd1a83544ff46751a777bbce23985669e43ff63fcdbac34d68f42de56},
  '{236, 1'b1, 384'h2c71abaf5b00000000fc949ada9b9b8923946346ef5af5650fb10dbee979f793371c30ad2f55ac70194b635702590bad, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hbc65644acb7dcf72bbf937e781d6de7bca052adcad474e3a2b06795a18db7b89d246a485d696b2b8d07c07d2ba2e2929, 384'haf811cb9772b4b3f1eed358b722a5b28a21617aea7eb6f9371b68a8d1eb7232def267ba56a6220f66a03c3ed7cd322e1},
  '{237, 1'b1, 384'he99162ce536e0000000093617fa47895f4b9723f71611138c0f5c75ab8da14e39bb777da07b169e146b4fd2af589752f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf6205c154a9cd38a1fc9a18c7bf6350699c95144268ba4ca182a5c8d50b780d468aa9beb8115f8ec489558891ecd6d65, 384'h863f41412ab418fe037fd688a9f6c509bc5535b2c6b5ad7bf9486fb0e5b02136219aca2cdd9d5d63f9140e6d1d054201},
  '{238, 1'b1, 384'hcc79f0ddaa267600000000adc5aad840e30d828999218f6601ae7a66b325cca1fed100d1c4d16be31ee15735bb9e9fb7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'haedf7382965359c9abff67f0fad2be6b84d760ac95da1c656989f19938b046371e101e8bab9a0ae9b9ad2bc242a98201, 384'h9175511515a01096b4d77cc505c60facfceb1841948442448e5c9f24204f817eb20d12479305e82ee5a34bd73ebb04ad},
  '{239, 1'b1, 384'hf201649bbff5243e00000000b075db6e9f524f148ae559a8d6892c2ff02310d5964db32afb47655c9917544aa7996954, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hbcc696d8d3445960e00c9f76f277e5fa3267224d0187ad120f9c074597eeafcb6c7f22f51900351848855b20072afdae, 384'h935dfc4f7b48ac01116e5cf194fd2feed3cb28e72cba8485f1d94e5d20f5f4147a1ca3d6496bbe915913d21c4f5afbaf},
  '{240, 1'b1, 384'heff457e7b98ddc6f410000000020323edb6928bb6ff781d3a067fe5296e693bec34236f0e5e33e4739fbae34268c03a0, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hc029e49048921647659a042eb533004ea3487f22a7f2c471c43a5a2326dd03ac24386242c05698194b5c6171f08bb7cc, 384'ha92ed5f2c736e27711384a131c464f73852a7dd167b27c63020040d8de991a390ad76627d597ccfebed809f2f7f57b26},
  '{241, 1'b1, 384'hc8bc15912f7da2f2d0d400000000c0439cdd632d268200760a4ac187d17ceea4718473e21385cc5105bbf541ceac944e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0f5e1771ba1957fe8794c23776832ea40ec4fda999186f6c365f4749f07893cb55e972658c2d3b39a7b485193ff1d719, 384'h3967983d1da9dcf0105ddc383f599539d4b32b1bb8dae1a6fe0afbc9bff1e0952a32f08d161b3979a60bb6e49b6c7d7a},
  '{242, 1'b1, 384'h3d8e42ab2348b2becb80cb00000000bce2a640c87bedcfd754e89fc5d9c7d66d405aa73fccc84addc96f19637be09d8d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0939874c2f67090a900ad7399df78c6005fc4673e23b155df7471b31debd2174fea94e00180ddc1a86609eda8830b449, 384'hc9d71934a7222e415a01692c7274e5097d580dfe74175dfc0055feddfb414c1ae857051ce12c0ff25d5372751456622a},
  '{243, 1'b1, 384'h50d9e34b483e1cadc1f206f700000000554047ca9be5c7a947d7e2c3a860dddf7709b34eb4600bc114f2dbe9f0916dee, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hc35b9eaa9a03a36ba52b7ab207ff48925a0188d288b1ed25d7de8bc203e8ef912a01891eab8f8e3a7d0a948a26d35ab1, 384'hcf04105208f10af61240da6073cc39278fdadc0578bf40bbd0b0f601ed791e041a90a09d7c423a83f6cd047d745c4f24},
  '{244, 1'b1, 384'h5b4e4b16787278c52da3da2b14000000009c2aba426bf6d9227e0e797efa1e0be4030776e2a64bcd4bdfe60580949d19, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6c1fffcc270c9bf108289b42514e57e3f29ea0f1b3fbfc10ea283b3e6d2a4438d591fb7274c9ffee15009cd9e340f106, 384'hde38043b47c7d5ab21d8ec5a35758f1a69ee59ea6df525884a04210172e7421f2a49f5921a4eac40b278f6e7c49474f4},
  '{245, 1'b1, 384'hfa1831e4a2112a431e6b9ba84200000000005c4e9a04d7169bf3a0be2ed8b063a9d3fa1f21672d2f5bd9f116235c49c6, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hecc637f3d32bc9a1ec20f025af72eb03df49f27901fef6b58d226b6eaa9faa6374f87c2aaaecd69946f3777fb9d4581e, 384'h48f6a06b296a17d84dd26ffded0c5dccf177e6df9a7710b0406fedfd269b2c220f11c1e02cea42c18ccac768c64ba7eb},
  '{246, 1'b1, 384'h3dd792dca8c7227014a578ebdb4b00000000319798a8d9e45b78b22cca7a41900db7c8b1bd01205e2e7856198a7c176e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7dcf9ded94532d50e9a2ac971642da0de95a1ca95500621174113c1d554f21bb2d175b5beacdd73443043c6cc8eaf105, 384'hd4da518de6b8c05c640a3e7a1540482d935c4dfdca7544daf94ac8135804127b93665e1191b66bdb0089c49802c33fb1},
  '{247, 1'b1, 384'h6de328a089eadf427c91e3da01618c00000000c874d1437727d9c7dec71ca6bf781bca4194cd94741f3f59ee4b8382ad, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8209054bb408eed6ab65f4bb76223d509ea24d02cbbc5273145bcb40189052540e565fbf50474f83db3da054a793c863, 384'hb8169b12568ffa03c0e37d4a19911e9f4af7cd256343a36e41cd7b41395524235e86d55c647f288fe5cef2b5401e4413},
  '{248, 1'b1, 384'h5be10e9f0a420564ff205f9817366d1d0000000000b298349541727f79b7a122c5a07749596b825d1539f84eb774ad63, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9fe969770d630bb938ca2282536f71f3dc461071186216d940eca10fc53c4e7ef067bca237bd6a82eafef0fb8d38050e, 384'hb23a042178fdea5da86229c08a51227f23e31b1e2345defa12ed7041bec31f87837ba4764721823ea9f1e652d536c5ed},
  '{249, 1'b1, 384'hc2469c63d410a38a627f18911e47b2ad00000000fb90d317d4cad91b84618a3f9b95c476bd91f1d881267b621125d19e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h459be510bca760f75aca10e41efb7ff64b78fb9711e72f224373b9af14f2c042b68b15bb189b3d7ccaed9318936543c9, 384'h579c07e99fc9891498ef3109360017052cb20bafb290ca2ffa64a72cf01e38e12770ba0ad5e190d2ef10c2d294e099a2},
  '{250, 1'b1, 384'h330a4faa9ad071616eafe267ce678db6ff000000007b042233297aed66d4f04ac127966cafd855673066fb4256687aef, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2bc3bb18191a5bfe6d13c735104d78dd947854cf1d93017695119c8f04ebb44d7a7fffe71d15b78e0c2c28765bbdfc38, 384'ha9051dd102b20e3c69a01a36b85a1ccea670da784038989145e3cd9108b064d6d54f7df21164adb91b3850cd005ff68d},
  '{251, 1'b1, 384'hc8d71b76b1be589043b9a170ef94f5087cb800000000ad41ac80d70a3f85ef372b64a927f0f40a6ca06930203f6c076a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfe2c0567483ecbc6086a24160200a9ce91e6cf52df6d25b2ab08fedcc4ca95cbb6be68b58870c10169264f3b3e8d552e, 384'h34b7ef7c580506d29b1ef8223e2131602dad9fbcbce6f846de42519faecfa612a82e999cbfed45f377b77ae5ef0b4835},
  '{252, 1'b1, 384'h1055a2316a22b80def10109152b84ed72f7c0b0000000042130eb1017c83d06e3dea36ddb2acd54f7478b6090b8ab790, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h09296917f12fb3bbe2c69c9bbbccf8a400d7e0b31c453ff7e928a7e4347a185435490790f56a5a819271192d64d612da, 384'h163860e1f6390c0ada261d2d0346b49f18ec3b17e0389e4c3b2296382bc23d6576bb968120cfd24ce735a14d3167f203},
  '{253, 1'b1, 384'h08dae202d4925b821cdfd4ff2fa8651a8490d50000000000984d20a1f372beb9186cc7284093fad4f39f6f4f6858a7bb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9bf980d1d91fa0daf73e3bcc02c7773503f291b3378c96700ecd71aed81fb8ff47d4baa8b6782842f227a9314f343e44, 384'h4342d335dd870f4a1b817b519ab184710c2c79b6329ae3f87b735e48874b6e47950db7c8f0fba59a349112bd2b3d9eba},
  '{254, 1'b1, 384'hbc9c5461f59dc6568661a5ef292204e6622cdeca00000000777d716ff0780d1137eda9773ce1ef25abe31e339c151ae2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3f9b09855b47d180d60fe6ac427458a452ad72678d13818d1a28a376b31fd7d1c67e70ec234c40fab7d17719f7caa27c, 384'hdc1d5765bc5c266a39e1a94085983ccc63cb41556e3733330c98934c329eb7e724e12cadd082da23952b831bcc197f18},
  '{255, 1'b1, 384'h1dbfea46c443eac946b540f32b644f021713502bdd00000000bb62e1d981bd904e1596b4deeddaa5c6c24b53cadaa728, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8c6910c012fb1a5b45032b09f2cfdbc7c3b22b0e18a0cc0ec4adc296cbfca66832379456b867ad1a0184ab1a80af59ee, 384'h3d87fec6feb833d01e4f77a306441fd27f328d01f6c20eef9b185ad4723c46f5d15e7be0db1c496018b4fa1987ac6b78},
  '{256, 1'b1, 384'hd7ab19e1f3b38b0e899222e078dbe179e1626d6b6ca200000000a8a255668245c6f348e73cc6fa7592de96d3a8a8335b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8cb0ad263557318156ffde6b45cb6ca8633c3b50b51454605dd01242dda44c9cc5b59b327e919629a9f73720e53a5e63, 384'h4f2a0cd11c7ac03425e25d84bb44149117903cc4638e2f64450e2a915b14c6d9c74f70c4f85d6036bc604a92f9b97166},
  '{257, 1'b1, 384'h4ccd1e431ee9f7555b25f8802ea9c2c07fad1e66e31588000000001ff77cf56aebacc79dbbccb4fc14006733b04485c2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h17d2c9d32253234b36a02e59f99163913a7c11a723f7122c521dba2cdec36bdcd1837c8b60a916aa64ed32b2c400d23a, 384'h821fb503cb89385bf9a6288ce6559cb69652e8bf940ccd0fa88aae2e72d31ac7d7cf51433ee45889094f51a4cc17272d},
  '{258, 1'b1, 384'hf6a91b683fd947e8bf0e6d449d1970fbb504f44d616d74da0000000095a265006c5371a8c74575faaa5e42a25e5b2749, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb2e6fbb2a70af41654fb5d632fcbf9dc8a8a362394e42d13e086e7da261aa980b49c4a610a367973f798b9aa9df6d0d1, 384'h6d237b3161ec602529eecb5c7c706020f82b8040ccf7082576e3caef5e8d6cd87c46a8f3ea9947b18d1a35c83494d849},
  '{259, 1'b1, 384'ha1aea299918ad61c922b29e972f8b4bb050443f573ce1ead6c0000000020c8f93a781adca4c049e601e9a3bcfca48632, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'ha6927125459e31afc31810117677c6ec2ba27c3ee5cc5fafbbd74153d3d2b2f7c7411e564c09d582dd2d5a201ec2b0fa, 384'h6e14a3955d24c4ac4f8c035f5edaf74e45ebd95a27954bb1c11fdb00fbc7156e96318d33725c0666006ae0573f7df785},
  '{260, 1'b1, 384'hfbf549b7f63be376a7947cd300baa17eff3ccc8d449cbf0a9fa5000000002ce01c050c896dbd80e886750a1b939c9977, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hd0f8e8a570a0462ea8ccb980789acbf243cbe946522ae4e9e6fa7e5e8e1bc006c8b84915355f00f39a61dbe77d2b4b9a, 384'h0f1ed97929bd7cd633f835086d2241a7b7d8f857b94f71e30b3e9bd19863a401834d01d29d32399006e8f84e0852e3d3},
  '{261, 1'b1, 384'h5331c588ac1d7a7f18ecf911e3285baaefaf6b504de84beca4bfd400000000d199828a434a003fb77d77922b6fac41ec, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h19e5a38c81ae167c70ef4a1879b7dba0dfaf5dc8a841269e82b106c6ea3f9e3f7e162b8c561d8f1b7b4a2cfba4c8a925, 384'h08c41e654d262ea6e1d2f74cd99ef479cb36476b2dac5bf0f250d87f7115bdcb59ddda54abf3b3b77471348facc0c8de},
  '{262, 1'b1, 384'hfd06f7859b95fc71f9ffbb8df32aabd3d2a882f26227863e0591cfea00000000c5b338026ff3ba3a1d5807ce8a2d4872, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he47a0dd0507717c29d0e482037d7fd001eff3b80013688085ae430d46edb23cab8df8716d078c6503e38a1cf6a9e74f2, 384'hedaf65e609db0925dff88d252791db4a008d9b46e5e6da98e23a766a8a35b8df79ec189d272429dd64ca60983462daef},
  '{263, 1'b1, 384'hc0caa5bef25fc10f618db2b4b8d2e3f7950505d21ea9dd312ad88c9f44000000001aef232fe1ec496fe841813061b544, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h35d47a723521553ea0440e6dea660439c51b80e896877b03b0c02ffabcecd86e6cfed2e4fcd80d76c97ef945b626b025, 384'hdd61311a4d0eb024288fae55abef6f0fdaf71a55cd3ccb2f8ba8d43ef36dd5562c07d2b4ef60e04ec4c696fcd052185e},
  '{264, 1'b1, 384'h328b2d7830d44a378c73b6da3de7a6d238baaa7bd85292556424843c884d0000000094e0f707b75177dadf65ce6372fe, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h5319f4a01c4e88261146de213d65e55c2532d9a535bc8c47cd940fd2b7b5bb363e1932bdacc9a196cde39368d86a14f5, 384'h8afea330d833a1f3310aafef6bc27b684838ef3e57ac7e36c02e0dbf9e33b934dc7afa7418aabc3e6b0841eff09bc470},
  '{265, 1'b1, 384'h590dee3efcef116007e32b5c50477e7dd075f4a02fd33d4bedf7e3498baa97000000006ec8444d2dd7c8ed66578d508d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h5c51106927cb275b54a7c90f6ba69902f1b1a19e2ac4b76b8d1e41b86f14ff32bbc66f07d4be610ccde84af4e1401181, 384'h551d9901408a4d9a1a85fa17de0c7bc49b15bccfae095247fc256a048582610b6ba87bd89dc98859dba2df76d77aff2e},
  '{266, 1'b1, 384'h609422c689ef615b2b0535bd8ec18b8cce65d197a1bdacab3f46ced79d1218ef000000009341f3e66a6d1681a7c547cb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he931ac049c0b7bd9060a58b0f78d8d0b60f57caf647fe6476802c9baae7e06062fe3d1a1f0c6345dc7c530db32cad843, 384'hb83867f656b9fea099ca0678bd62f2013238bbd6969a2384e0cb2488dad615a4d91dbdf7908426c9ea9ecf17b872a25e},
  '{267, 1'b1, 384'h9b1af634930bb603b45145a699391fbc262c3c2945f16d310669edff29aacccca7000000009edf5c285270cda2b39bb7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hd4ccc6e89e85ffcca4b9e32fd45c5be1585d20c35ec83253f3080b0705746f0f5e7e92043b5ae8fd95963e45b4199213, 384'h48448f45ad0fc8d20fd1dbd088bdf6d51577f79a1e5e55432ea79d84eefe0b9b55ba145d637be5a686477fe00e1fb481},
  '{268, 1'b1, 384'ha900ee181319e7a92ee017d61f168c4266765e9c3e33ef32a9edf055bbfbb96949d6000000008c3bf70bd017a758b48b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6d3ea919365f9f39fe1f9b8c17415766f4c2b77c8393dc8cef321af5b4aa955646643ac32b2220b7590deadec15b88af, 384'h4d64a4fb9e26aaeec0d92270becbb5e2f04d812b2bb8b86cb1744437e62e58dc72f98ecafeadae69aef3328953143490},
  '{269, 1'b1, 384'hcfadd7ce8a12f10af606f03c05830e0a7969849a80924b77b31d4b1825ecd6c3d6bcb700000000b2713dd7084c2ffc6a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7774080a80e32087c8e923c65522c76648205d9804805bdf05977c4559eeacc518560920e55f626748ae12034745f7bc, 384'h1bfbb5bcaff2b70298456fd8145bbcc6d150d9f2c3d91d6ed0f3d7eacc16456f698138ab34a546195941a68d7e92f3be},
  '{270, 1'b1, 384'h5fcf143a3798aab86b588f5d30db580c5126f1b58d8a17d8154f01fdcd5c8d967c7045d2000000000c85eb6584638edf, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb8232417c371ecc56ef6342abecfa42afe479ad1cfcb18f8945ab0e2076621c185c2821a8028c36f1f2a8d3be7fc3442, 384'h17a0f7c15403a3fba3d8f095cd7eea597df761dc46e5c8122a3fffabb9fe37c52232e7f49af7e7cbaad8ed62dee8a371},
  '{271, 1'b1, 384'h3816985a4eefc2f0eedf0cf5cd65796bc9074daed0165ed1a36a1b96116a794823c8316e5100000000d9bbd2cfa57d6a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9a5e7ac2a195f5859a0753087da0a2ac20a8bacc551d4c19b10fffe6b7acdd3ca6543957c9f7be8bedd33e89df7ba594, 384'h106cb9821f8aadaf7a7c411df6ca3bde9b6d4a267e4a43ffa9d5d29cc973f3ca4d776351b82586be7d6e2c251726b3ec},
  '{272, 1'b1, 384'h70f42d203bdb579a69f3cef0929487f7816593692484cec51ca5f1caac122348ce7eaea2a849000000001a55c02ef8fa, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1cdc96cc7892322075399aac7e0a86d4ffdb6e45153c0afa98bfd912941c22d05f360fba6f8734542eb55375b26d38aa, 384'h8ec452f8acbbef3ebbff11e6bf349032b610e87946a6221cccb5055c18d1f1188b6254a60113ed8adc6d0b09fb2f3fd4},
  '{273, 1'b1, 384'h10aeed5349bf090fdf3f3987bf954d059aee8faa79a12ec6f845918992d30af7b51d20be06ca4800000000ed135a15a3, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h937d4df90d09299bd32bf354e1121a311a77ba0274e7b847804a40d5b72ecb8e9e441afc5289e0337ca1195a4951c1e9, 384'h7e442371b9991905f417e4e67ead31621bc068964097a46d5bda507a804f5b3bb142ff66d07012549fc42cec38754d11},
  '{274, 1'b1, 384'hea79b63b9dc825d5b1f06225f080e1b5df6aea661373d98ca5c6e0529a245bec7025be22acfc534800000000222534c8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h65210ed179af3b99c09b9e95dc81f77007a32002ee7d53eed567086a68a62f1c08543c85f7d1e1f081bae477ff3613fa, 384'h025ce6efa2fe24732fe11f5b1f1232d48fa5dbcfbd62f96776302b1ac52f0d0d40549f2b2f67299569cd14fb7ead4c45},
  '{275, 1'b1, 384'hb7280b7558119ae9a6ab3a9e950b5ff2de0142fb86baa1165a2ac5a1542e832241c28385ae8dd53f1d00000000506ebb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he6a4518771467967e264a9b736aa1f8bc6f421de607fec7e93fc62d91082c979930e6a3ffdcc54d5f0f4b4a2f0665d49, 384'h4c6c625b60ab3230e6d190f37a6f14e574f8dc7595467fe89ce62d6d1f2fd198368769fc84b556a3847be26841351408},
  '{276, 1'b1, 384'h1fc79921cffd33565750256ee48f4afe5097716fd012c1b64c1abfc96ceceade4ee8b967a50d580191b3000000000677, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6388afc6cae9421ba6c52a640a0ebcb9c547505f500307194c8c1eb41cac959686ffa7b3a2adda65136030cba17d1695, 384'hcb1e148645580dea5a87c60db7c818942d55f169fc59eda9a2177a001ecc1bcbf2d519d67d79fba44daa2945bd380c52},
  '{277, 1'b1, 384'h54532c36b250773519e5c8c0b6bbe5d8653b6c9550c439017998bfc1198b66fc5e664cfe7b454a909c52b00000000057, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2d7f29f767ba2f21619347bf29494a318eee949e91181ed7d2cf61162b92f0747c308885891b1734e9b6d5d3705475a9, 384'h1c34c2ce61e3dca2bb3202b6c4320155f764fc58d318ba44df9a7c06a0a453ee43b633353dbcfe129a54ddc8b6a27e13},
  '{278, 1'b1, 384'hc08b51e60826c23eeeac7be3cb937a3a4e9569f67811e2f2f0c701184dad0edc7fc31ce21c705040378b922300000000, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h68a8758fb66c0ee50309490852f214f6bd09dd888f35390163defa70647202983ebabff3791287d016164c945494edf9, 384'h099a2c1073815916cebd4a41448e1b8dc9bb150465adf99c8a965b5fb327bb879e1b34f8d7c509aa1b018f98c9e13e40},
  '{279, 1'b1, 384'hffffffff65e6a7dc05cc02c53a50a75250d0531a889967be08ed9c1cebaaf411685adebf5d765590c71698a98760864a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7ff134c055bda5bba91fa53da5ff90c501a6264abd8db5ced03e9eb88ee63325f267a8fe483b0f7f129434d2e2114705, 384'h11649294f067d415681ca6cf6245b0beadcb4095b8e9c9d18bf11ebae41ecafde7529796286ec2efa9073de2f9025e3d},
  '{280, 1'b1, 384'hffffffffff119a65525c432a989ad477745e7aa11c0e53765ec2ae6126c5a03d3e68732df8de98620f972a6420225b7c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9dfc836f6a993e1aeba9fe4b4e09901b83a5439a0ede150ab583c217fc22154050eb9c4a2f1f0f75c06139549d3013ee, 384'hed83ee554777a5086ac90b9654f724507a54e5651b4d38153ac7576cf8dc9487be7d3efca544ff4b4804981efbda10d7},
  '{281, 1'b1, 384'h6affffffff5071ff7c18bab2e95953b4f00b0a3b6e4f6d87ce17271f82688b9f6d455b89cbfebadc2185858abcd54d8b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfd614924d6325daf270efbff4db11d645ec9b1f903fd36e1543bbd536ee010d07dd154fdc945a57f52f239439279f42f, 384'h079edf2f7ab361f7542bfd9175dd41ec137bc00d997943720e164e7187585a487a1893cde536b1dc52cdc0baa1fc2183},
  '{282, 1'b1, 384'hd8c5ffffffff73816d056266092bbca055147ea761dd6d1cc84bd71cfdd5dc17686f9d30862585c8ff2a122ee3f23965, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'heb55101d2d489c0151d991b0e486016222997b917363f8c48386683091297819662ccc34381d5e5ec1c0c43d137232e0, 384'hd8bd992c2e0ab4fe46a4b43dc3b5103c123ca38e88e3c555385a6fc8ece7d9c957776667f389a950bca4b2ad6503c48b},
  '{283, 1'b1, 384'h8280c8ffffffff347c8fcd28a68e495ca9137a15e21c11291389fa92ff4a1e458dfba63ca7b442d33fabbc6b479edc31, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf29aea476f19eacc44749f6057d39c6da903ba5c5b5667694145a6fe053ee08abed1d6869d3830036a29b063b295e67f, 384'h2decfc3e7d8cf0391f8e21714eeef04fa4f660a404294bcab6cdf23e4fa9e44997694781c49f4539a8d5b0dfa55603f1},
  '{284, 1'b1, 384'hde2a1aa9ffffffffbd2071c366f0eed18d345eeff7644d11fa09bfe9220610aedf60598a560c50f1d4b42e9702ac2102, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h4b55c6c5f0264ddd31b88a92072d3a8f33b28306716d5430c0ff8fbc37d9ddf1e4a60e4e496b355f77ed005b51e352be, 384'h54d6da5a6385fa10e97c21b5bdb732a9a9c0685883da74f1f8dea0ae497b7609b3aa4ee92f448144ea2c5529ec2fc016},
  '{285, 1'b1, 384'h5ee333cb21fffffffffed2c55e54b05c5072e23b0e9df2ed91556d8a0772a36ce570fc4dc899a5f4adb6364c375c235a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6024ed7ee8ef3edc593a9d07856b9aa78972ff33b82608c93e7068bcac05e0c5048889c8d520351047fa80f050abf83a, 384'h0d221dba3ef2d3c14923a651bd2b803603fbc94634033d52a66d80ea6120976c8fadc7274d05ccd47e1d06a63310b6c6},
  '{286, 1'b1, 384'hd6436d5df1deffffffffd88bb9f4e47eec31ab00857bfb9ecf90ea403e9a65d6af9835ce6e2c1a77b870b719724320d5, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfab3f2cf338bd7bf46dada597a4f66cbeb336393e4a289e21f8a02a6428bcd5fe66e87bdd3b5072997f94b76f04d9aa6, 384'had0c0f1d9c4f8a4b5100e183dee6d5d6825296784cb8205d448204237f5d3435f4c8f0a4fef81890c5a5a028405330da},
  '{287, 1'b1, 384'h59bfb0e85daef0ffffffffc5c3dbc4d40b827bc0a1da0557c0db95cb14079a5e4e98e119c269a452a86fea807dc7ac1e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h15cd4339b568212b20856d8397e5c5aebf3b4e4eafd8c90adc2dfe93f928e8a8bf17ec307064ba866491d4b44440d116, 384'hba9357237d9d6b22be6761f63d91a265d1dc08cc693ae14576200d6aa7322eca439eea414634f5666c22ab29c67fbcdb},
  '{288, 1'b1, 384'h7b40e2bf0fd54a19ffffffff4c6f54cb9b82b6a7d62de54af61fe36d81f80af65d7f058aad786911e25a26f9012642ac, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9d2deb753b8e16e6f24e1b718000daa0d4617242225f1b91192b1ea8acdca607b05f1c0da8e3cdbdc52f448a376f13b1, 384'h8654d2738725423c0934c20b28327f7a5ac53a61f296a5ce562c8684d2f3090d19811fe70dbce71f106c4060740981ec},
  '{289, 1'b1, 384'h2f792de69c2acb0d7effffffff48117939bcd7d48fc75d87bed984c081057fd5b27ea9e2b46362c505a00d4663e1e9a1, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1c7c8d1c493bdb1f1290f04aed3c4a7cb0a83c36330a4fab50e68f235777579dd06a073a3857f226dae511a2569e928d, 384'h14e5058d70b7cfb04cfb0c3c1d3d6fe500328340860e4b7cc2b5f11cab09cba0c7b887274453ab30d9164c73fc1f6f36},
  '{290, 1'b1, 384'hd7cb0d5b3da1856dc731fffffffffeaf9aa058e75ebc0284acd14f28673787a2fc2b42c5538eaf5031b96fd403d3b0f4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcade486e6a8e78141b15dbe60095e42d8196fafd843c722c8c686a60063e701f30d8a488c2a18a63635a13bc8ff0a787, 384'hed7aa0208952d2d452432ffa1bbf7146080911cf7e87aa848ee90314b2afe427a80cd70187b3ac3572a360d4db6b17e5},
  '{291, 1'b1, 384'hfac48e2f7fc095232aaf2fffffffff54095545e463574aae8f4f277fe0b0c1b79d5e1bff50b6e9f07b9883ee6e2818f7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2787240e7fd6d895098d1773733727ee5792fe644b0774b8530ddd758b347143d1939bb7c9a3312774cf7126e499f5ab, 384'had215cb6681f287ffb96a6e7c41331a2e773e68791391c658f2e5c95cf82e3871e49c9fff08f7b540848c1a7cee2ab85},
  '{292, 1'b1, 384'h0e0104d1b5eec3d01aa30c46ffffffff011932f39144bd30bc9bb51d57dcf4e5d6a7ebdd12cded759e97c62016e89c1c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'haa92d0b7d6046210024b962fd79d1a27ee69c25936e5895cd92224b3f560829c11de20e7f52320bba91b87c4c7ef4962, 384'h816c95ee54c677c4be1ba70317a90aaf1c1d2f233fd480d22cab453d9539657ce695e21952e6157ce3460680dc2fdbf2},
  '{293, 1'b1, 384'h5b045006f1acbf669f78a23737ffffffff4a6d9156a79d3842a71ea5dcdb3d1591b682821e9397086d0788698a7c7ab3, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h4eda9fc1e0df8ef24f3148f8a737a76eceddfa6057441c877816ac402349f32571c8074611179968e6fe7cfc1f41a80b, 384'he0549e78e774377dffb9e742f05f5b1a1a2198571d0f2243fd25703029e0effac2808fad1c82efbdf0063d6032df33dc},
  '{294, 1'b1, 384'ha0282563c4b28930a556425c4e66ffffffffa8e5ad6e3a31f7c0d0887b2467b179f6948cc41ec8b3f1317956536de7d4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h18a83b96dbd10de3a62fdab7142f201f9f480447bf000f6ee314da64d2351bbc7bb94cd1c551dee4828a603e6a853fca, 384'h8fbf2a1a7ad4ed76a08748f41f5b3468a9a7cda57503aa71c455292bde2dc88a2580a65a6859d20f924aa7a5cea3743d},
  '{295, 1'b1, 384'h79f16206acc319a5197163434c1e78ffffffffb50c8e19d5fa72c72b48f5ba71c64a9386dfaec75aa3c82368b41a6c9d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2fb5726226521d1105cdd22e84ff46a36768ee4d71e6f5cfe720ddbd36ad645c05a7207c9f7cae2d8236d965ff64f943, 384'hac3f8b7841b31c95f27e99a86413b6aa9086fcdbd176f7de65a696d76edcb0775f2e257db75fa5aa716946f3d80b1cea},
  '{296, 1'b1, 384'hc000b06ba2beedc670436cf7b895472fffffffffeab748f165633a1585bbcd0d0b91965aff1b0e9627a6dffd363743c7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2a38f4cc1da426f15d8c8dbed58608eec86862554f4d6d503dc6e162e72754b1298ad4508ae2a93d493c836b19548c4c, 384'h9b51610514136d5dcfda3c4736a839288bc1f043ea362cf6e56dce3f4337204d5bdf92160a034f459b30410872dbeb0d},
  '{297, 1'b1, 384'hda248a16e5573a906c85cbf5e8ff6ea512ffffffff37e31bf41b94670c215f394095ed5c3dca3767c180bd8562aef90c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3407844641a75ba72ed05f9b7289ea2c8f9015c97e8d7aacec4a88b374a255371b19e7a2e7949f4b78b63334b4984434, 384'hcee117c6fb8f8e47ce33357d7ed1a82b1ed912be3778eda9de303b2ee910c014eee3cf03e27f16fd94d7ed5a8e8c7b05},
  '{298, 1'b1, 384'h322fc62ca75b7741ac679bed13fe0e4a782fffffffff3f459548e73678d16fc987bd4e505188b3f2121c65b5cdccc039, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb98e1313e62ff0155158059e422cb6e8ce70d103f1a95a77e1795ef2ae38a42596732405602299ee730b81e948083adf, 384'h8a34134e86354d26f343343c05cdb46350b610ad16883f234e847fad97047ee4b8dfecd0bf77479b65643f9c35b74441},
  '{299, 1'b1, 384'hfb9a8f07c555acbddca310f455bf11263f3488ffffffff5a491c4069cff6c54a5805efe17fcbb76d2e1fde16fe7ac746, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0ae0a9cbd0de42e6590835374548708df9671208ab72e23bf7aa4329bbd0d4a696e99d04d36534e895737b468cff08ea, 384'h8c8b6bb101ee844bc75cd2b3b32ea9c3b6c2ac5408c26f6a444335d730af2dce6f4bf1bf4585428e902f901eed10da62},
  '{300, 1'b1, 384'h02aa6fb89f1d295921cf5564ebe3b40665ea06c5ffffffff7759f3fb122187bd4509ae8f919e0bd2a897b8299d07b9cb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcf0310487690de93d344bba957a1ba380f72c2ae44975f69716b2aa2a866787dfc46629825ef19e5528395d872ff9367, 384'hff60a995865b6f5e6ffc15884e5901d55f384ffc62982e54a9c2dccaf7543246673c5bfe710f2a29daca77de766ee9ee},
  '{301, 1'b1, 384'h286843bc06e8c45270197afdadbc2b3e0622f8deabffffffff545f876be899d7835542fc303ffa3d6f00e14c5ae2a1a1, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h4a0f3d91ef6b9b6e512cd9c996f8e896717ea8c6d685834e4c31bcaf592a93d0f0b169efeb0ea52a5bea6be361d7a7b3, 384'hc3d429d0daf1ee7c2bf4a0bc8f10cd7ce453b8e2a762b31885d36f5e03cdae3adb693bc2efe8a64d6e7bbc17f23b5500},
  '{302, 1'b1, 384'h0c1a555d6e050dca35cc8393a58097ebd1b206c335c7ffffffff8465c1af66a0524307c757df1c8f2e5d902d44e6652f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h40f82935328e34e31f1966bd0bc1dfc2adf1d71d86fc6dd0f9e9e1930dfc357e30fa67722c562dd84cdb73fb715b622d, 384'hcf40658591f34527587b0969a45ca5a30f87dbcf0b058f75c158ac883d52119030881c0aeb1f8e12682d06d072705550},
  '{303, 1'b1, 384'h5d331817df8aea58e841ea2b7d430ea4d7d3dfddfcd354ffffffff3f98e2f7bd1af8c469965458f0bbf379d73a72b1ca, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'ha3434df3d065f4b32957077f429bccdaa8875981006ce880585c160fca1f552dc6334583d7698226e650e95d86a896b7, 384'h54e2eb28c70796e3bea9f2fdc3799f7d6dde5b3cc84de7448296d65fd8a44260b0666cefa416adda5046f45a5b8a9ae7},
  '{304, 1'b1, 384'hc9954b68f1638653fcb8a41e23d6dcc020789b8cae823ad1fffffffff493db702e2e33241c076d1ef7876411c8bd24c7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb54b004489e12ec91e875f3062dff1f1bd0407e216162b4913a34f19943c8f967c1f7250ff0ce5f43a0b250bb9fae16b, 384'h95c13a702ca6269ed8cac69291e01767c0f862648b0961238ef0b6be88cd316973a290bae4f50147816a49ab014a7d69},
  '{305, 1'b1, 384'h4154b64bfe35bcecbee1092972ab973511cd26e999d8beae7dffffffff5f6a3552355a24fe170e7ae4cef52c97da7996, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hea28a6b9158328d0711bfd10019643648e695c1fa9df2a7c2e1a6d3b03b6703bc763f8f0c701d7b925d35075da783f38, 384'hb4bb6b034288af213ecabdcc2d55610181ba77b26673b1490e7e08a43f6e57fe20618a5adc7fbfcbe255fa79655aaeb1},
  '{306, 1'b1, 384'hee00ecc8c6860c71fac74e858cedb957432ff7f8489a47efa6ebffffffff6b75e29edd887bb98674f3aaa39b0d8ddb1c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hd973f5fa26a7069dac82790097db0d93dfc52a490ac2a84960c6dc52c2e84d2df1917c8d194789fe8981be40fbefb006, 384'h1dc1ab55752add3952ee3f5d86bb167ed1fdf20e19d5c893c1a6031c1a2b70701ba03cf7d78b89331d524c5dcf38462a},
  '{307, 1'b1, 384'h8c863fa4d1107a42e4fdf154ccb85f80f45faffa10d9ab2f0f3c9affffffff87671314227064df4f548b7938a98547d1, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3d4ed5e71127a0da4aa63cc1d7ce517a450370dff65ef95b4185a44199181ec5ff70f80f6d7435e6bec4d6e58e73591b, 384'h27b2d65bf08ab8e745544225181638af5df08b85c9f7a9057e1605f145b3a1389661d9c990d0f4d82636dc6332b6941d},
  '{308, 1'b1, 384'hf09c119db64dfd9324626ccd1d982e02d602d085ffbc4457a3d52effffffffff288c6ec6e9a545a1ae9431eae26ab6b0, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he36ffc2ca7e62c2fe35c7761a78ae2839d1503b437cc7a89eee28ec74d75d2948c7a3148070ad715f7ce8260c160611d, 384'h0c18edef913d63ac220cd4b28aef1cd43aa9acf7b0fe889c4a28ac22934e46aa2a99a5b803a61471bd5bfeef8c86b17b},
  '{309, 1'b1, 384'h59d5aa030e5773e64f85e1480d80e1137c9e66d3a78460dc051a4addffffffff08bc0d6358eaaf7b236dae6128f23dba, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h148906bcfc686aa3f608321d17a425373bd9ce2f47a35a6a01124992cba56e744daef2b00dececff63ed96d5d7c2e158, 384'h4303a5c7049766956679f204e655301dc16fe9cd85f6ebb1997410e0d2029240181c946d86800cc6ba882f276603db29},
  '{310, 1'b1, 384'h6a88dce7f07d6d241d8ff668cad03e95a16b52d89911663972a1bdf97fffffffff9577890e6980fa4f66b10cb5d6b8fc, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h5264c26ceb0481b74472f26ecca4459785a2d63c9494d8744e42e9eea5799bfb0fa95ff3c8a5de2868098a025110bbe9, 384'he1858d96c814dbd39ca5dbde824be0894b4e418fe51306784a8fd0680850a5b32958714ae9124e9ad6372412212df1be},
  '{311, 1'b1, 384'hce8f67e22a3012b0a74cc986fd0dce36552a4b3a3b6664c575a26de406daffffffffdfe12b3d8a4af5358647b44249dd, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h273e229dddfaa7ba5763c8563f3a05c7d2d2471331225e8f26a20e0ae656115c62ddfac3895f10012253ba7bb79a65ca, 384'h89a6ab6fd5bca31659278ac3f3e79ded9a47a6fd166fc746b79fc3bd9d21e5f332bb1e89a14efcd3647f94aff9715aba},
  '{312, 1'b1, 384'h40c6210cec4684dca0928c5d5738f6bdc588df3d78f78888d21e0a7ea72b8fffffffffdbd60dbbd4720725d0f7c0f495, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf447dcc8ce6573a2da5fd58a3974f46a8d76608e477742b68c2e93245f359567a953cd18dc1d95fa7e3c5d02210cfc0e, 384'hb273a9ce5a021a66f6a44f2ae94f2f5fab6e3b5016648c9df38756a5b7e71d07aa453240d39bef0d22afab1e19095694},
  '{313, 1'b1, 384'h6246fd756393fdf4b4975a5b23dce0d026c7135feb6356e4050cab2cd769d48dffffffff95b1f61223666a16e8660a3f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9378874a38f221b27d8b7ab06d827130d0db2e9c43f443e9cdd254ef77a4f7aae589a6c1499970dd5acf516802688aa6, 384'hf94a6319379598119bddf9f787e74b135ad193b692e44a848ac6d1d0443d49adcdcf1a9f530686e76080840e1b647be2},
  '{314, 1'b1, 384'he0968793bac4ef008e53ed3760a0f35b8785bdaa1df7f2650234239a45bcb4bd75fffffffffc4ac022449381ad1ef3df, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'ha48cc74a1d39a0b8cfcd12768277535389790c9ad2638aca42401a44e80ff0ceb40e193cd9e27e39443a1d2665de485c, 384'h1569ca82e563df78feb1d704953b8c35b7eda09259fc16ab262304d0c09383f550cfdc97ce549874212e3fc7b83f6d4b},
  '{315, 1'b1, 384'hfc16b96a1dcc08d5f4dbc5aa9b1d7ba93e0a13bde11b4cddfc429d5278648790cb2cffffffff0c081b428b25d09c041d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he6049a43aa5761ad4193a739da84c734f39f2f79f8d97241982082185fe9cef7747b68c59ef3909f18af6c5df48ee559, 384'hbb7800436791bae910fbfc6b69c0b7e6972dea1bd5ad82aaf97ebb85d920a15f9f5f280fd813281f36b2ae3c53fd6e41},
  '{316, 1'b1, 384'hb61712846f6ac1bfcdc1337eb9d69ce264d6703b585dd60f2b59869299a15afabd6ab0ffffffff98662c144a2e76cab5, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h148d734104a52c9d58ca1ad7ba56fd35147e8d324a0923ebc9c5d8b393f492bce1da6c9d1fa68d4faeebf0868e03f171, 384'h4629809043f228f0f3adfc0696c2e9d800791ee82034c5fac37fc521e40f9bf2250c53036b8286e032959ed5f3a58483},
  '{317, 1'b1, 384'hb23bdc0ab0199b13e19fcf7a9a65897de4f7a806c84ec41fc99fd42a86f30334639d4db1ffffffff9c2c4ce9990579ac, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h16762ba4645c905590e6a3dd4b1e2af693cc4e64153812f93b80ed4d1c07e664e5b22880f24a120d4b48e1400fcd3afb, 384'hd481c2f9b255bba2ac29fe055536c3c7fa92e4f34cfdc5b5f5227f582736c87c1350bcb760069c4004ac33fbe2ed3549},
  '{318, 1'b1, 384'hb72a59d0ecfda2bb05e0ae8d4e0ba8265044b76174980887d64404d98b9aaa26b9500159d1ffffffff220cbf1a43db70, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h830c8c92465fc7f1a654d22eaeadf62b5fa29bebc8e184ca104913eb8bea234d287961900f308d88f9bb7387c8de58b2, 384'h960eb635db967cd69f80123e0a43501c6161cbd9e8058f5bb7506cc24fba3a3694688b5b0e066bf2ccaecbb5a9eb0c9d},
  '{319, 1'b1, 384'h74c0181efbc542cd0a9eb39d63ad27282ecc3c0d0ec4ac94e5cd96fa60d54856bfc5bb34f4b0ffffffffa87f077fc767, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1377906f42629010e79bc60142234a44c78e8887f6dc4086bdc7e9bf94c92c84aaf48efb0269205b8bd6e324224df178, 384'h6f430a1937fc0463143c80a0e132074a64acc825c2f4ed8b0de03204a681bf171e9e002a88431fd388c7a906511171a4},
  '{320, 1'b1, 384'h64f9579e23ebf443e57d6a269eda73e343b673dc34cc55a14d276ab7a73c2bf244dd4cc17e5573ffffffffbe3989e7cd, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hd1d335dca83a7ef4770e68ff82d2bb75341abf72a362c88d8a176020db37bfd5874e14c0cb011cb316bc6e6d1322a893, 384'hc61fc7dd9f66b8cf2f8c9a780089fe31a20608b458ea12a246a1cba34566c2d833a71bbe09482ad3c26bf9bb6088fd5a},
  '{321, 1'b1, 384'hcdee4a1b6555fe2f2de30ef0e9355f08f24640183d29d82d8fd45b0953449d481ff5ad9e28994554ffffffff98e4f4fb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h536183374fa37f210723fe3aabde18997be247be006e20c5d17d8e4c79790ddfe4e6f17f8823d36aceeea22c9e44ba9d, 384'hb6a0f63b27876d1686b9e601c273c20530c765e506605cea39d9accba9a7007bb10d64333e5e22125f34d1dfc8e60461},
  '{322, 1'b1, 384'h34d149372065fadc240fb01f2b5743ed462c3b2436472e74a69d3feb01f4600a051c2cfb1fa51a24d4ffffffffde2b23, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2fa6073fd290a699ff0a4bd425a69d4e151a3ec3faa65c504d5e41b45c2a738d343a99865690bcc22c03230c3949ce3f, 384'h3989dd2d632007c498ed830d277cc1193590f23fe5e778deeffdbb2c135258327b121a81313a0bcc9f77db206afddd8f},
  '{323, 1'b1, 384'h326b5d0c7aedc94ed25a2757b94cf4f6d28a23e4b9643f5e69b16d952ba6875e2e054b4b7f3ea63fc09effffffff8f82, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcf60fb9789b449ac9b9f022dc83481777675e55f09b4cba5d8349c0e16907f8929e3b538cce4d71c01b010a633807997, 384'h67654a0bebf3a63fa93cf9906c846cf5edbb03968c86eef5e7555a14d606009006f9f9e4569be3375a9a8aa04aa20c45},
  '{324, 1'b1, 384'hdd29193b789fc54b4f2494bb4a077638302270d27bd7b66555f7dd1657d6cddafd31433fb385ef8b5a2affffffffff0a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6ab23c76784d003ec508233f7f5e6461d6806c66af62c4769d45ec8751d276bdb68b2efc4fcf83f675a3101941f9adec, 384'h6f306bd6f782aba3c7d0c0d6c0e0e8897f967f0de2a84db1d67e477378ea425dcc6fc6113e5a5f67ac34eca2c69d0bdf},
  '{325, 1'b1, 384'h66bbdf6b95d0db8ec971af150c99a68316ac3d07e92540590a73e0e3270b81eb745595a686d480f58fc2faffffffff0e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h526365e36472883664eb011bdf9a1503397f0e3509066665f9c276e367cf2730774d4525125cadccfef0c0cf28949a2b, 384'h948cbaf1c0e7f0ccca5f5d2a7e4a94f4a7ec43d2cf69ae5ebecb41521daa9e618615208cb62b35809fc40401670ae3b5},
  '{326, 1'b1, 384'h6692e0535e44ef3757292e65849818d0855787f780513f5c82d4b1ce4101510cd5656a20dc213c05cb338f4cffffffff, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb1cf39b023502a1aa3daca372c295c1eb3c5fee2a841ef2cfd4087ffdd4e35e8804b8d879a939216d24fae1bd1e7f19a, 384'h8b8bea55a9625efb9733d1dcfad8d426b81c9e71fb53b246ae54c3196972d284172e6b1911bafe6b631e5e48344c4409},
  '{327, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hd7dea8ac1e4b9aea2d3d1ad7d6a877e116a8bcdb87c8463c69ad78f8074f33b2c179ac0580af901d21851cf15b3a5e34, 384'h2a088198c090b9e367695a1c7fa110b66828d8f07bafe6eb2521dd20e517cebd295cc9cce52e0c0081b4cf7fe5ea884e, 384'h000000000000000000000000000000000000000000000000389cb27e0bc8d21fa7e5f24cb74f58851313e696333ad68b, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52970},
  '{328, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hd7dea8ac1e4b9aea2d3d1ad7d6a877e116a8bcdb87c8463c69ad78f8074f33b2c179ac0580af901d21851cf15b3a5e34, 384'h2a088198c090b9e367695a1c7fa110b66828d8f07bafe6eb2521dd20e517cebd295cc9cce52e0c0081b4cf7fe5ea884e, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000fffffffe, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52970},
  '{329, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hcba0cc097c795cd467d835977764b7740fa480c3cad83a726d68bbfe8dbb752934eb4fb6c767dc09bdda6d0d2d057ae8, 384'he277c7ad56d6f21099d998e7bfded8c8d2d100c8ebd9f57681a633b91ad0890c020e724689c6b1b4b8f35b49679a4fa3, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52971},
  '{330, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hffc271e311cefc1c133202448e2ee74457bb68951b0e575747cc6ee9c0691720bcf9eba23c18f96e845cda05e06d4f7b, 384'hdc7c5d17e91f12abf3638fc8e87866f0373f0ffa90c2c759712d3fb163730a184e4707ef424ef833079c0ed5e1498344, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hd1aee55fdc2a716ba2fabcb57020b72e539bf05c7902f98e105bf83d4cc10c2a159a3cf7e01d749d2205f4da6bd8fcf1},
  '{331, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h74ae987af3a0ebd9f9a4f57be2d7d1c079c9ec7928a1da8c38ff0c2b9bd9822fa7603decc1becabd3f6ceebb353cb798, 384'he0c9ac6f4f575fa1ed2daf36224d09aa569f8b1d25b62fbaeddf766a34b9309000cce2447017a5cd8a3ce76dd5428ff1, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hb6b681dc484f4f020fd3f7e626d88edc6ded1b382ef3e143d60887b51394260832d4d8f2ef70458f9fa90e38c2e19e4f},
  '{332, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hdc23280ae627109b86d60be0e70cec0582a5b318fa8254dfcb97045eefdf1aa272937de99c6b3972c4cd108b4fc681cc, 384'h0ec5438a5d44908c479da428e5b2e4f5ae93bf82b427d8dca996e23d930700082828112faac7f710928daa670b7576cb, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{333, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h9bdf0a7793d0375a896a7f3084d3c45f8dfcd7f73d045484e71128713cab49b4c218af17e048fa6dbe32f2e289ee8395, 384'h0be28a090c2f6769f85e5ff1cfb300bd0ae907b5d5367ede98dfd3e6a81c4b4903289973285a4ef91b790ad12761321c, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002},
  '{334, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h90770515f27351111e56d3bf14fe392d42186cb870374a8d40870830057bf52da8c2e27691236a0de2876893f9b77ab2, 384'hfb1cb5dcfd30e3a2a0056a5dbbc1c5d626ba669cbbfe8bdb121de7cc394a61721d5c3c73a3f5dea9388cad7fbca72649, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003},
  '{335, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h90770515f27351111e56d3bf14fe392d42186cb870374a8d40870830057bf52da8c2e27691236a0de2876893f9b77ab2, 384'hfb1cb5dcfd30e3a2a0056a5dbbc1c5d626ba669cbbfe8bdb121de7cc394a61721d5c3c73a3f5dea9388cad7fbca72649, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52975, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003},
  '{336, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hf7f5f9382da5dd3d41cc2d4e62570b581b67dc2ad456de3af75ad1ce7be27af8a77771e67a08f2dc87ac91c5a744886c, 384'hf7194e819162862cb7c39e39445da63adfe10704ef7407f1fcef062c8f86729c700da4f9e747c5c77e32dd25e7f867af, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accd7fffa},
  '{337, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h24f0d59e6bab85cce63823e4b075c91520e0f7090c58dbae24774ef25917cf9fab1030513f4a10b84c59df529bc1d3b1, 384'h2469f23a674bf49a0383d239ca15676704eab86bd3149ea041a274643866643b786bb17c5d0f10dbf2bfc775c7087cc1, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100, 384'h489122448912244891224489122448912244891224489122347ce79bc437f4d071aaa92c7d6c882ae8734dc18cb0d553},
  '{338, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h39833aec7515dacd9546bab8dc740417f14d200bd26041bbf43266a8644628da82dbf53097fe43dca1c92b09832466ec, 384'h67f862c02c8911343a146fddc8246c168376e4166e32bad39db5be2b74e58410b4e9cc4701dd0b97ba544142e66d7715, 384'h00000000000000000000000000000000000000000000000000000000000000000000000000000000002d9b4d347952cd, 384'hce751512561b6f57c75342848a3ff98ccf9c3f0219b6b68d00449e6c971a85d2e2ce73554b59219d54d2083b46327351},
  '{339, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h6cc5f5640d396de25e6b81331c1d4feba418319f984d8a1e179da59739d0d40971585e7c02d68c9a62d426ca59128e0f, 384'hfeab57963b965302cffe9645cf3ee449846381d82d5814e8ca77167ccf4c20ec54278e874f834725d22e82b910c24c2a, 384'h00000000000000000000000000000000000000000000000000000000000000000000001033e67e37b32b445580bf4efb, 384'h2ad52ad52ad52ad52ad52ad52ad52ad52ad52ad52ad52ad5215c51b320e460542f9cc38968ccdf4263684004eb79a452},
  '{340, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h567e0986a89e4a51ff44efdf924e9970cbdaf5796dea617f93e6e513f73cb529e7a666bd4338465c90ddd3f61823d618, 384'h5b252f20921f66a72dfcd4d1e323aa05487abb16c797820f349daa04724f6a0e81423ddf74fdb17f0801d635d7af213d, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100, 384'h77a172dfe37a2c53f0b92ab60f0a8f085f49dbfd930719d6f9e587ea68ae57cb49cd35a88cf8c6acec02f057a3807a5b},
  '{341, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h95512f92e55b5d18003397b822c1173f4e25a2640a4a68bb880a6ca8605cbfb83c75dbddc4937ed822e56acde8f47c73, 384'h48e4ff027a1b0a2d5790f68c69923f3231ac61074caad2a022f6eabf8c258bdb8142be43ffa16a6f2c52f33cba006400, 384'h0000000000000000000000000000000000000000000000000000000000000000000000062522bbd3ecbe7c39e93e7c24, 384'h77a172dfe37a2c53f0b92ab60f0a8f085f49dbfd930719d6f9e587ea68ae57cb49cd35a88cf8c6acec02f057a3807a5b},
  '{342, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h74d5679e10edc41eb06ba54a1de2c9c71820bbac14f3758bb7fb593dddbb2e573e0d7a785344961399da18c8f615ae1d, 384'hf71e1c0ea892931571da09432ac46f6cbf53129e1e3e74c567180c037df59da84c8374b295b5a0ec6100ce9d800cd05e, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc528f3, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{343, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h1764c83ff4c28f7b690ca1c4b05832d78394f0aa48de452eb7b470526f4099d45de563b506c1570eb9b0f899a5f03f5a, 384'hff89e562385d77b2c5d48dbb54501960997566bca5dcdee15848b907ee7457f8e46a221f64091c36f8d3053147c1a628, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{344, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h1764c83ff4c28f7b690ca1c4b05832d78394f0aa48de452eb7b470526f4099d45de563b506c1570eb9b0f899a5f03f5a, 384'hff89e562385d77b2c5d48dbb54501960997566bca5dcdee15848b907ee7457f8e46a221f64091c36f8d3053147c1a628, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{345, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h100fd7ac4ae442ab989f94a10a1f310f799d76980d00a14418db067b144bf45fa7639446fad508b76fd3ad9c9fe55810, 384'h693598529b8349a28dd1d0632039ff0897523fed9af2356c0e36612135ed629369448b97d165ae5b2fe5c5ad396d2b06, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{346, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hd9a08d4f9f8708471e2e6b04ce08750c395b80f4a14169123e2fd97556c1171d82e87165a77b2dfd089ad25382ef4251, 384'h517d0c26bebfce8483bfb089243d82eb0e712a7d2e7f71f9abb82ddf16c2e525146c7dc5686fb7ad334022ad092d32a4, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9},
  '{347, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h68133653284ee7e9a8cccf584a9e4f06bc31a3eb031999f0229db7c2b10630424c7ee7513e40319e3972c1a5152d5d28, 384'ha547a17df730d86278de44cc099643ebe1f07e48618de255bc672dff63c58f86b2db29c89f109147d8d6be1f03c466e5, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294ba},
  '{348, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h233c399596e090c132c8e8b33c2ed443d73ab9abafaece5e47c6a6dc82d3fcc006ebf8b5b1c5fd028c97097909d5be38, 384'h035f777dffaac0ef909bbe6be4e01ecfae3b36b2ea2095e352c179737980f96124d45b76677274d975eda57436f453de, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c},
  '{349, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h357931297f6a369df1e1835ae66a97229c2ab63a75a55a9db2cdbf2e8582c7c0d8aa79f2c337e4e01980d7d84fd79917, 384'h06b1de385965ae26fc38ab2b18a8ea60e52faea5c2e27666913858917cb1cf5b5c0bdc9c1498389c1db155e54d3198e2, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h078dcf7c421b705191d0c45a27c93d16ab513eecfcf7c9042fd744d6d8dcefe1036fde07248d32fcb19c725c0580a027},
  '{350, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hb760dcee338ca73c8cc69f0360d87253ef3632d302bdbf743a65f8762ecea207a5c5aff3add177378e133378d2c83a40, 384'habcba73c686f35e13d1cb44197bd763b5221d3b17ca7d888bbbc52eb2c33462036dd7a3b569290cb586d9e6514d69b92, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{351, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hfa8f96db8c7c9350d90ab49baaa941a79ebe62f017d54b6f83854f430408926e4a46335e44e1d67f0f18c7db2d70ca93, 384'hb65df386caa193875fe91740214526a2ed17393d8bb62bdcee9f887802bc2d76ca9a304b94e795032956c8608c0e7f46, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'haaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa84ecde56a2cf73ea3abc092185cb1a51f34810f1ddd8c64d},
  '{352, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h69bf123fb0d38b6a1c3f01a811e16ac78f40301332a0a18454fb4bd9b7c9516520f5ace9eddad328b8d283162eed1c75, 384'h9fa36f89c13419404c11c2ac982777cd30aea7e621351d96ba39676c26b36ccd109035d708da63ab9aefee3c82f6d405, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h52d0bad694a1853a24ba6937481240f8718f95b10102bcfe87d95839091e14aa1c38ba8e616126d4be6fe25a426c2dc4},
  '{353, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h1e5863f2dafa6a4d1a10a4cb18ebe792c0154aced0c5c2abe33f727335c720693e92749795539350d8503f209da1bea5, 384'h6f0889c25cd0aee834431262177f43b7ddb01a75532dd55086c44c1931cdd3e0312eea51d300050130f6e754aa9f92f8, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h2412cc835da0a4357d1b7a986a76fe42b79542258c02dd7af927b27a9f9352ed3eedb6520a422e876949cb5fd0724090},
  '{354, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h87fc8357860b94528775f3787406b79d7a7d65d23d1d5707e66978be71aabae87bc539c24addf6c55468cea11cfb85bf, 384'h3f881573285dd3742ecf062d5321c3d5f86212ba88ae75dd3945ebb3b44c37a178d440bfd72ca8f2e7c99cf6367da248, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h1a2303bd73ab20717627366a498a23f4afe23f30b93b0f3be65b74e5eb19f2abef049411ba50146a305c5bb98169c597},
  '{355, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'heebe3763025894619173c8b4397deb7febbfe10fe2d283fd303d48691ebc8ba3ab1209278e763199a18f398b9c148405, 384'h98640539d7ec66d3c43bfed723292c85856f02e020deff4e468bf3bf3c7fd08391d9525a2cb4f85fbebbb7945a5853ad, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h2805e063d315ae83078dcf7c421b705191d0c45a27c93d16a277765a9f34e9a4b2e3bac6291d3ba508e5769fdbc4920b},
  '{356, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h41a0504da3995adb7665654b6ef7d0d00f77fcc536fc1cad41b0daca5a60dd88c99c20e698c99d5663eb532a57db08b3, 384'h4d2b0acb79b95b70cb0a5e2eba110061ef87f0d34b5bbfdeaf5184b67103f8a2bdcd20a7b9f09ad11811776659becb75, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h5e063d315ae83078dcf7c421b705191d0c45a27c93d16ab4ff23e510c4a79cd1fa8a24dc1a179d3e092a72bc5c391080},
  '{357, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h45c152c4e642f156b50ef6252f2b0cdd36f20cfacbe389fd79e2fbf19f0810cfbfe5d157d2fcc9b2a649e9675fd86c07, 384'h4eeaab3bec18eff3b702e0e0f5c40ce928ae48161e06833ef3d76fa743c51b2711ca7c06cfc3a20ab804066251d2a115, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hbc0c7a62b5d060f1b9ef88436e0a323a188b44f927a2d569fe47ca21894f39a3f51449b8342f3a7c1254e578b8722100},
  '{358, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h5f6849efa9aafd6a4030018579e39d241df4c192e5ba78c6e9b441aabdac8eb8f4b353865c1c9127ecccca468c41a561, 384'hec501582456fe6396643c368d2b9735c47384dbdcf2cc16927ab9b327c36350fe7e1f949e7ce14e60b1c1dbec8dff5f0, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hd315ae83078dcf7c421b705191d0c45a27c93d16ab513eecce49d6742e48c5aa2b36ea79df9d9e3277247c3d843d5887},
  '{359, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hc3ecd74e383f55b7ec8cf0579e6fedb9863ee0a82cc84cf13854dc1017aecb2a5969f15194a9ccb09e823559fcd7b6f1, 384'h1faa3cd553119de6efd237b9a84dfe520694ba373c8b60d5b2e741b35bbdd9cfa635353a1f0cf47042881684a96fe516, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'he2c087faeed9abb45e3942a10187bd6d2df94757e2584ca7599b3385119bc57f7573f71dfcc9161dd86a91096695d236},
  '{360, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'he4efcd7525aa87a1390ca91cd3f0ad38613384377278c4e29b14264ca550e6e57e6c6559df830065caf902a2f8df41ad, 384'hff1121276e4228ac454d62994ca1a3cd24d500a90ddaaee2e5203da658504292bd81b62c4024a8fd4d0725e6a07c254a, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'he727c7f2d36924d4f4fb46d5d0c752e8aabb5317b2e59419d1d54ca40b148e12b60908edf846b56e4d64224fb8d7e885},
  '{361, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h54a018053bf8dff69ce32e1f8c0c9ba658dffcfc1200cbd89c16996aece05b84ba945164b4bcdb4d8b6dac967ac78c47, 384'hedaafea84b25520478e67b328def37e5bdb94f18f3bce507cc24161aa4297477fff23968ae367cf0c3f2f70ed2bc205d, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'had2f45296b5e7ac5db4596c8b7edbf078e706a4efefd43013f89f548eb1919353be15323e74f80a62e7c37108a58fbaf},
  '{362, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h68828912c312ed14280c954102f2d4ab06d58bd9e7abd0afcafa0c349d0f09100bc5c91156cefeb9d3e33721f5d1d5f4, 384'h69cc3a91967d5b964963044ea966e4a3e2488f3be4232f1a8723d2956c687240fb2f92d456bea0b087b1007b444141a9, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h83c6e7be210db828c8e8622d13e49e8b55a89f767e7be481fb9d492c668a0ee02dc4f5dcb69eed3bcf4445e36922e4cd},
  '{363, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h1dc3d0da27139b88b61893d1bdee2e5fce3dcd8c4b65e1861ad0886068d32d905d343c4567ab20903f43beb1f5e3059a, 384'h3cb44b0793c790e3f65bf78799755a8f40107cae627b57fbc03181f65b12416ba5f5fed566a95dc4b1b93a1a63550811, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h8d1181deb9d59038bb139b3524c511fa57f11f985c9d879dd6df6133efa89045a38f50e201805df28ea43a9227177785},
  '{364, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h85d1e93894969ef05e85263e3751285abf14ce1fb1a947d99ab869e61249ab515224ab3b0f322be36c90a3a1522f83ab, 384'h88fcdd8457e34a9e8105d361fb3711b544e4684aac178a3217505bb894e851181033d7c756d572abcea1aa7bb1e10c6e, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffed2119d5fc12649fc808af3b6d9037d3a44eb32399970dd0},
  '{365, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h609b7164d1e196a5596bef71b34a8fb4eacbbea10fd41d126c16ea3578d893e898c413805230c7fd7e33ee832be72120, 384'hc2e379c857c01d95b53daf382fa5c196705c7f927ab3dcd8e6aa6bd4fe6767c56c178dcc1bbde32ea00afdc1a4f59fa6, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h79b95c013b0472de04d8faeec3b779c39fe729ea84fb554cd091c7178c2f054eabbc62c3e1cfbac2c2e69d7aa45d9072},
  '{366, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h6f557ef52d480ea476d4e6bb8eb4c5a959eacf2ee66613dc784fff1660f246a1765e916d20ac0dbc4543303294772d12, 384'hdaba49f78c8a65d8946aab0a806140136516cff6725267865e9f93e4052e072ae984f3e975e7792b67b5b1807160d429, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hbfd40d0caa4d9d42381f3d72a25683f52b03a1ed96fb72d03f08dcb9a8bc8f23c1a459deab03bcd39396c0d1e9053c81},
  '{367, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hf07a94c4b1dd878c2b4507549ad7557cf70f7286b95d7b7b48a0491a635379c0032d21d3fbb289bb5b7214e2372d88ee, 384'h38934125ec56253ef4b841373aea5451b6e55b7e8e999922980c0508dc4ffd5df70627c30a2026afbf99ef318e445c78, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h4c7d219db9af94ce7fffffffffffffffffffffffffffffffef15cf1058c8d8ba1e634c4122db95ec1facd4bb13ebf09a},
  '{368, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h61f352564999c69ce86c0336c9a9a9baddcf4555b675183ea27f682a7b0661250ff7d2d00672880e7d3fd5329b4d19a3, 384'h1f28c529832d0b336633e3ef2b0bf97007a61b7e427c9d2ca1fc2910b0cc685d409ec423bf2f5211742b8d3b33d2f04a, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hd219db9af94ce7ffffffffffffffffffffffffffffffffffd189bdb6d9ef7be8504ca374756ea5b8f15e44067d209b9b},
  '{369, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hd23d62e8f8c286da7a8e2aaaad9b759c6852da31639ebddf7b4e4fd1ebe26806caef21c9fdccced05cbe1332bce4bd4d, 384'h899480daf03c5918b474d9dac0742ed97aa622d18b747c4446191b5639abc708c02ff97147b5092cc1395da611476001, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'ha433b735f299cfffffffffffffffffffffffffffffffffffdbb02debbfa7c9f1487f3936a22ca3f6f5d06ea22d7c0dc3},
  '{370, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hd1c1d5980bb20f6622b35b87f020a53d73fe7d148178df52a91964b541311bd88e00b35834238a0bc1401f9c3ea0c3e3, 384'ha50b861b701099048e0b36ec57b724b781f5c9e9d38eb345dd77eab0cb58b4fdea44e358bc6a6ae4d17476eb444bc61c, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hb9af94ce7fffffffffffffffffffffffffffffffffffffffd6efeefc876c9f23217b443c80637ef939e911219f96c179},
  '{371, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h6626339de05be6e5b2e15c47253ad621ae13fd4d5de4e4a038eb2127fe33fd5b898cd059a43ec09d186fbf24ed8c00d1, 384'h9251db17bc71d07b53e8d094c61b8e3049e040da95a885e4e476a445f7bfc3705f8c66a7f7d95f0697b9bf2eff9e4cc0, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'ha276276276276276276276276276276276276276276276273d7228d4f84b769be0fd57b97e4c1ebcae9a5f635e80e9df},
  '{372, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h6288739deb45130ee9d84c5d7a74a64d4e1a829a657c8f06a178438b8657169c486fe7c2610ea1a01b90731edf8e2dd8, 384'h1f2d7a092ecf4a08e381473f70519befd79e3b1484076fb837a9ef8065d05f62df4753a26f72162f8be10d5bdf52a9e7, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h73333333333333333333333333333333333333333333333316e4d9f42d4eca22df403a0c578b86f0a9a93fe89995c7ed},
  '{373, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2bdc91e87927364f316799ffabbfcda6fd15572255b08deb46090cd2ea351c911366b3c55383892cc6b8dd500a2cbaef, 384'h9ffd06e925b733f3f017c92136a6cd096ad6d512866c52fecafc3b2d43a0d62ef1f8709d9bb5d29f595f6dbe3599ad3e, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffda4233abf824c93f90115e76db206fa7489d6647332e1ba3},
  '{374, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h9aaa6c4c26e55fdece622d4e1b8454a7e4be9470e2e9ecd67479f2b7bb79ac9e28ba363b206ce7af5932a154980c1612, 384'hcb930ccefbd759befafdb234f72e4f58e0ce770991dac7c25bc3e4c7c0765fcf1dacbc55f4430520db7bf7da401080e1, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h3fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294bb},
  '{375, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h9004b1043628506e37308dd0107ba02d809b1504f89948161ab7a580b9e2b6c111688f9a7db9ec1e52c987cbe06f1173, 384'hf20b953d46c6172a883fb614c788bf860c456b1b08db110b09447ef0176f7222be4120128f8a198f37264efe6256af93, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hdfea06865526cea11c0f9eb9512b41fa9581d0f6cb7db9680336151dce79de818cdf33c879da322740416d1e5ae532fa},
  '{376, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h23c5694ec8556343eaf8e7076de0c810ce26aa96fce9da325a813c4b0462553d679c70a3d9d626deac3160373bf05d11, 384'hf4e0f85a87d3b08a699d6e83d0c8309e7e1646625f7caa73bed83e78b2e28d8384f2c0555bd1023701c10a2c1726a9dc, 384'hb37699e0d518a4d370dbdaaaea3788850fa03f8186d1f78fdfbae6540aa670b31c8ada0fff3e737bd69520560fe0ce60, 384'h7cd374eebe35c25ce67aa38baafef7f6e470c9ec311a0bc81636f71b31b09a1c3860f70b53e285eab64133570bd7574f},
  '{377, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h23c5694ec8556343eaf8e7076de0c810ce26aa96fce9da325a813c4b0462553d679c70a3d9d626deac3160373bf05d11, 384'h0b1f07a5782c4f759662917c2f37cf6181e9b99da083558c4127c1874d1d727b7b0d3fa9a42efdc8fe3ef5d4e8d95623, 384'hb37699e0d518a4d370dbdaaaea3788850fa03f8186d1f78fdfbae6540aa670b31c8ada0fff3e737bd69520560fe0ce60, 384'h7cd374eebe35c25ce67aa38baafef7f6e470c9ec311a0bc81636f71b31b09a1c3860f70b53e285eab64133570bd7574f},
  '{378, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h916e5351bd3efecf755786fa77f6acfecf3b00cd496fbcdecd8d255120dfcf27b70e7fc9de74be9b15f72650b3eedfdd, 384'h5bb6bcbdf478e15f77221d01d6086eae7dae44a16bdeb4afe178eb444600452789889310ad61014a3957436a59a3239a, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{379, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'he79f9ee594e711ae1439a237a0db174abd0b0138c4da3db1a6bc0180280b83020104580528d1030544ee4e7a17341e5c, 384'h393de20f319b72e523b0b9ff9cd10cdc4a5b6b35850be57079e1afd30dbd6d4651139cfe0b16b32b074f81563009f7d9, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h33333333333333333333333333333333333333333333333327e0a919fda4a2c644d202bd41bcee4bc8fc05155c276eb0},  // OUT_OF_RANGE r_len=49 s_len=48
  '{380, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h9d91680bd5ac912ddecc5b609094a8d5fd12b5d5af7c5bbff8f129d9bcedd5dea45df2d09513ec7aead188885fd278bc, 384'hd968fbaba2bd7d866f6853a6d79661fd53f252ea936573f6bc7a32426c6a379d3d8c1a6b1e1a1aa7faa7ffdf5c4b0fbd, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h33333333333333333333333333333333333333333333333327e0a919fda4a2c644d202bd41bcee4bc8fc05155c276eb0},
  '{381, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h66c48ea217602f3e0e77f402dfd386450c3a33f3b9a266d01cfa4d8cb9d58f19e7cc56315a5717ae27f931a8b6401aed, 384'h0f47cc979e0edb9b7970ac66bc66315d3d38594dc933dfb963ccd5676efb57b14be806c0879b3cd28fe6ddeaaaf4ad92, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{382, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'ha03d026431e0f75a9ce6cd459eb268c44d59a00bb6facd5b816a2823845e7f65c48c69cfb4841bc0ab8c981e6c491db2, 384'h488eb2d9321b30ebf3f1f99da618d3311b01928ae9b23764b530e2ad41dd121b6812b7a8a80f669934dd8efb0445a962, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{383, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hdb12e7908092c195819ea7652a2f923f678f00aa8181f3c2cb0021e268a176737d48a48ea25a48ea2b0cce3c31f1406c, 384'h9c46a9b415ca03d1b309c5f4735b6ce48da4d32a0eab51772dc6bb7e63d835ea7612c92a629c058af638a5bb5354110e, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h6666666666666666666666666666666666666666666666664fc15233fb49458c89a4057a8379dc9791f80a2ab84edd61},
  '{384, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h532b95507ca92950613dcffe7740715af07953e881d133b75989426f9aea6ed1bd22a9eb899441b29882a8e4f53f1db2, 384'h65dda7154f92c561b2b6c9f154af3a589871f5290114a457896fd1e9af235de9f1eb7cfe0911e27cecaa30f90bec73b4, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h99999999999999999999999999999999999999999999999977a1fb4df8ede852ce760837c536cae35af40f4014764c12},
  '{385, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h1dd1d7b6b2f677d7e10fa14bb35a74bcf83d6ea0bb308ffeb7d73634f6911e4213752173fa76b2c5be12d752b8176659, 384'h888325cc90b23ae34fac03a5b9a30cbcb9d24e02923d6d68e8e54066eabbf8a87272827fb2f26392dc45664bb2399e90, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'hdb6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6aae76701acc1950894a89e068772d8b281eef136f8a8fef5},
  '{386, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hedc6ddb4a76167f8f7db96dbbbd87b241a2477e60ef21f22d0fb235fdd987adb15a13a9c9f05228ec7e33e39b56baf17, 384'h8397074f1f3b7e1d97a35d135760ff5175da027f521ee1d705b2f03e083536acfef9a9c57efe7655095631c611700542, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h0eb10e5ab95f2f26a40700b1300fb8c3e754d5c453d9384ecce1daa38135a48a0a96c24efc2a76d00bde1d7aeedf7f6a},
  '{387, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hfebf3b365df31548a5295cda6d7cff00f8ce15b4aa7dc8affe9c573decea9f7b75b64234e2d5da599bf2d1e416a75007, 384'h69205229d1898c7db1d53a6bd11079458cc40da83c16f070e5772b1d2059fef19f0f36d4471ad85ec86cf1cd4e7d90c4, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{388, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h8373e65ac625a5a4110e350e7f08a0392f8261581c06a88b125a145681687fc5a6c796f16ca48977bbfc7729bba80063, 384'h01d966a2d30fdf2b6dbcc8c9ac3b6b2150431f95fdf49e8ea5fff99f185cbcd2f9631ee3f074d680700fe693b0398583, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{389, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'hd8b5b751bef246a3769682966232b714b05d99a37199223e55cbc4df6941b2529e57965c94f60d88837cfd952d151abf, 384'h9eb51727dc4665f8e74e8f5c79d34ffd11c9eab8b5b773950d1f2c446d84c158aef8bbf93b986d9b374f722d94f59f1b, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h6666666666666666666666666666666666666666666666664fc15233fb49458c89a4057a8379dc9791f80a2ab84edd61},
  '{390, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h5f2098bc0eda6a7748fb7d95d5838a66d3f33ae4138767a7d3e221269d5b359b6456043b7a0973cf635e7424aaf1907d, 384'hb1e767233b18988d95e00bbb2dafbb69f92dcc01e5cb8da0c262cb52924af7976d9ded1d5fe60394035cc5509f45865c, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h99999999999999999999999999999999999999999999999977a1fb4df8ede852ce760837c536cae35af40f4014764c12},
  '{391, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h018cb64da6154801677d34be71e75883f912274036029bb3cf2d5679bca22c9ff10d717e4d9c370d058ddd3f6d38beb2, 384'h5bc92d39b9be3fce5ebc38956044af21220aac3150bd899256e30344cf7caa6820666005ed965d8dc3e678412f39adda, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'hdb6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6aae76701acc1950894a89e068772d8b281eef136f8a8fef5},
  '{392, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'haedfc5ce97b01b6201936777b3d01fe19ecee98bfade49ec5936accac3b02ee90bd5af667a233c60c14dac619f110a7a, 384'hd9b99c30856ef47a57800ea6935e63c0c2dd7ac01dd5c0224231c68ff4b7918ef23f26195467e1d6e1a2767d73817f69, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h0eb10e5ab95f2f26a40700b1300fb8c3e754d5c453d9384ecce1daa38135a48a0a96c24efc2a76d00bde1d7aeedf7f6a},
  '{393, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h3617de4a96262c6f5d9e98bf9292dc29f8f41dbd289a147ce9da3113b5f0b8c00a60b1ce1d7e819d7a431d7c90ea0e5f, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{394, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h3617de4a96262c6f5d9e98bf9292dc29f8f41dbd289a147ce9da3113b5f0b8c00a60b1ce1d7e819d7a431d7c90ea0e5f, 384'h078dcf7c421b705191d0c45a27c93d16ab513eecfcf7c9042fd744d6d8dcefe1036fde07248d32fcb19c725c0580a027, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{395, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'hc9e821b569d9d390a26167406d6d23d6070be242d765eb831625ceec4a0f473ef59f4e30e2817e6285bce2846f15f1a0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{396, 1'b0, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'hc9e821b569d9d390a26167406d6d23d6070be242d765eb831625ceec4a0f473ef59f4e30e2817e6285bce2846f15f1a0, 384'h078dcf7c421b705191d0c45a27c93d16ab513eecfcf7c9042fd744d6d8dcefe1036fde07248d32fcb19c725c0580a027, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{397, 1'b1, 384'h0c63a75b845e4f7d01107d852e4c2485c51a50aaaa94fc61995e71bbee983a2ac3713831264adb47fb6bd1e058d5f004, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h9da5c054a9eddabf4753559edd5a862cdf57adc0c2717a6949a43d80cfccd02b14ec06113ccf08081be43552391cfb16, 384'h88bb307e9a04f923c70013db3ca716d21b313dde0cd6849435bf3b192d5266589a00b34e9c4c626b1055e7a38ef10853},
  '{398, 1'b1, 384'h7e8809d33f8613073e25a0ab5df02a92dcd4362133c25ba5ec3d938d462eab421d82360a9f7969c2435e564df636600e, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h22b0ee0e8ce866c48a4400dd8522dd91bd7a13cc8a55f2814123564d039b1d1e3a7df010688dab94878f88a1e34a905e, 384'hf7668925262da6aad96712f817a9397b79f0fb893aedcd7221f454a60a18abb3b165aae979f29d22cfab18fb61945f87},
  '{399, 1'b1, 384'hf8723083bde48fae6e2f3ba5d836c2e954aec113030836fb978c08ab1b5a3dfe54aa2fab2423747e3b4fa70ec744894c, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h3db6c4d7d482fdb0a13470845f5ad2438198776c2a5954b233e24230889f3023ff64e4cbc793c4e3e94318b4e65f8cdb, 384'h03c22aa010ea7247ae7cc6c7d0f6af76f76ef91ce33a028de49979bdc2cc17d7df4c19c0e4c61c49275bc408697e7846},
  '{400, 1'b1, 384'h4800b6ae1095611eed9f358c814f4a35811a36349fecdb25c028e77019015896cc5b8ef1135d359fe1e24e8f546e8482, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h7a36e2c2ebf9bc0165ff75f5906a4806c2a668cb48477f7f105169c9b5a756abcc06b05b4d5ac42ecfd12cdd0f8fc65e, 384'h96aff9db7873cd2f6aa85c2693e1129b7896340287762854062df8104162a4572bdcbaf673af28a92314ec597f7acfe3},
  '{401, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 384'hacbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'h82b41176571a051a82c18e1ffbf4f3ef7146e0634755ba30fc965efec684d12830ed366acf4759fcce146e867b9108ea, 384'h52eaa43df5a95a92aee5f0002f4b4a1c870cdec040c966280be579a15e865bebc1269b084e17e727bae14b8ad6e6c73d},
  '{402, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 384'hacbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'hb4c1897895e4c214af7ac546230ab6ea733a6353fa11bd5d9892dc89e113dffb50a3581e58d5cac31efee0d56601bc84, 384'hb1494f4cc17f4baa96aa2c3da9db004f64256c1f28aefd299085e29fe5399517a35ae8e049ec436e7fe1b2743f2a90a0},
  '{403, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 384'hacbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'hc9b58945eed8b9949bd3e78c8920e0210289c1029cdb22df780b66aee80dca40e0e9142fc6db2269adbc4cb89a425f09, 384'hd672273cc979c16b3336428a60a3627bf752f9d7f1ba03c5e155cec8fcf523376feab08fe0e768f174828adcd17da0b2},
  '{404, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hd1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 384'hc6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h9ad0ec81fe78e7433ccfe8d429ffd8cc3792a7ed239104ade9b7c828332a5be57493346c9a4e944eec914acac1ab5a45, 384'hcab9be172e51ff52c70176648c6c6285630594330d8ffa5d28a47a1b8e58ec5c32c70769ed28bc553330c9a7e674da8a},
  '{405, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hd1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 384'hc6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h84ba925242eaedb53cc529e4763d8995aa7315e68a47ef89f291dd29ef138e4810bc1c58a6bcbada3ac83541dc139c79, 384'h4579278b73adadb63599028b873bf5f7cee2ff01eaf0faf2d529b01211a63e78433011da37fab174607fe90a4c3d81bf},
  '{406, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hd1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 384'hc6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h56a69cb5b4026268e11631f7fc35830e8a612ed79278f280e7d7e409558c43ef226ab25cf639aae7f435545cc4d8e8e5, 384'h5066494754680d61c23419273ba030df0f0b8b0a486cb0dd498298a34db478a6c133b4f5e071b6696cdbec63a74d84c2},
  '{407, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 384'he6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 384'h6328e30a8e218904631d6e8858e1e3841a2f6c0959af1b53ad3515bee16cbb600b5abaa5123c8eeb8cdc9b2da1a8ef39, 384'h40e708de5a00178926cdb263afcb12710ae8c03b298eeadbc40522c0479a94e98dfbdce493fcf0cf7f4afb6949d9f95d},
  '{408, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 384'he6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 384'h34b9ce48ad0aac78ff138881f3b13badae7e1cf5da7ff060c5642b22c5ec4c76fd4cd46d564676d4631bd567a7ea9284, 384'h61dae7993b4500005f45f55924c502f8803455e21a62499db2cbbc80a582c1107c8014afb4619f5d4d37fddbdf2d7bb9},
  '{409, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 384'he6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 384'he337217405a8457b0e31ae4e909eabe79343331c4dd0623c2b13d0981012e28d1fbf88f0101c1abae8cace1c801dfe16, 384'h948603710e13fe5b87e96ca87fb17bddb5762b9e4f2fc6e1c4acf4ee20b641518158b32bbd42884bffad25e0171a3462},
  '{410, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'h000000002b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 384'hd1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'hb2f22aeb025c40f695850ca8d9243d671557ecdb28ba78ad2f3389e78fe685251a29dfbc2ebc1d7e5e1098b4b286db18, 384'hd2ac24a65d1463405bd4bb117e4d1ed7f7d9b457d51dcb1fd8704ad27de5cbc11bea45f8e3cd1ecdb51981962feaa4b6},
  '{411, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'h000000002b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 384'hd1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'hf3b374deaa912309be3a08722fcd0fa17fbad8a0d674a96b1140efe2f9451e373029546b84a565dd88b6816b03c69912, 384'hf44fcc8e2513a2574e9c88de1960e8d7f6c607fb0aa6400362ccacf86e56cc44bfa6e233a993800fe1385e747312393b},
  '{412, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'h000000002b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 384'hd1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'hde778636b0c8775a48e8f7c2da3ce056ea18c0f7b61a6ceebccdc1db0462a739a9f623b342d82b5cdba9329fd32d4870, 384'h5f843dc49e8c8642d0ade1fbd635ee1ea6f6da8f980ec1d839de2b37ba7082668179cb80e7c97775e77c7afe8dfb9791},
  '{413, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'h00000000208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 384'h8f6f35102ebc10571603d65d14d45e2658e36a961d790348df0ed3ee615d55919e1c31d02e48b4c29b724e75094e88e1, 384'h1674424d64d3a780b031e928ee3b246a3703868aef1afcc6b50dd217ae6bdcb5fc7f59d2b14dc4dd08f22853abef621b},
  '{414, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'h00000000208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 384'h81fdae0b7e18cca48e0bae1a4e2c96f3973b0f661ccae269c1f0535265954e76473f51710fd2eca0b014e0386bdb387e, 384'hb4fd60411ae7ad836c8b1768bf44fe126d753781628a2b34f21fe1fbc961d21a153d3838e0200ddf8b7c16819230c0e2},
  '{415, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'h00000000208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 384'hf6b94cdc2083d5c6b4908063033dbe1817f5187a80fbf21e0155ebc16c3b14b06282171a63d8c6ad173bad8aa40b8406, 384'h569db82936c0d284c752149034a28e2415b57247c723077d8a5a7c9725ebca7603de5b7a41c53fed2bed8143a9bb8beb},
  '{416, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'hffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 384'h89d3d1a5c2ce6b637cc9e30a734ea63d34a7a72630400ee82916b79fa9a9a83b4e2faf765ddcf1fa596a4c026293ea06, 384'h9013c5c51bde3c114ae0ce19141c6c72bbf0a8f75885257f202240af212064f0fa9b1409d8c5e195a8db9d996eb1cd67},
  '{417, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'hffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 384'h4bb0ddb7af2d58e75b17f7ea81c618ca191efaa374026901fc1914b97b44ed64873404b40c249ee652e9685c67347881, 384'haf0bc80678b411ce0ea78c57f50bbb9b11678e001d92f2f49ad17af4759c7a013d27668ed17b13bc01e13eb9ee68040f},
  '{418, 1'b1, 384'hcfc55cb4b6f445aca0641b0ed200bbdedef9351f80ee5090d8d1a90f45cf2696786caa2d4fafab455b15678bc517f0d4, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'hffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 384'h024deac92bccdf77a3fe019fb5d35063c9ad9374bf1e7508218b25776815eb95f51c8c253f88991c3073c67ca8bbd577, 384'h8da6b6f9fde42f24536413f8c2d3506171c742b6a0883de116b314d559388b41630aa24c485e090fee5f340c79486164}
};
`endif // WYCHERPROOF_SECP384R1_SHA3384_SV
