`ifndef WYCHERPROOF_SECP160R1_SHA256_SV
`define WYCHERPROOF_SECP160R1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp160r1_sha256;

localparam int TEST_VECTORS_SECP160R1_SHA256_NUM = 70;

ecdsa_vector_secp160r1_sha256 test_vectors_secp160r1_sha256 [] = '{
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'hc0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 0, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=0b(0B), s=160b(20B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'hc0d64c9119a1ef31b0b0b1422b8186ace88a078e, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h3f29b36ee65e10ce4f4f4ebdd47e79531775f872, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{241, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h2a08a7f52a3506c5ff0b0bdfc41ed256a998deca, 160'h3d5324b851f80f334befa39b77241cf06535a1f6},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{242, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h48dbbef868af35b058bd34e507e85fc61fd60f31, 160'h2efb7e448ba59de5835198c3d5f5015113a3dae5},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{244, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h47398e906863d57ea273977083d36ce35f1f619e, 160'h24959c9b1f06bb8822bd8fac8f45945fd1c7ebeb},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{246, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h4b24155af66bc983050381c2579ad91a85c48d4f, 160'h28b0d445e93fa372a59b7030c67d2124b9bbd65f},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{247, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h57999b6dcf7d77337d8445543f1ee0d212d7f85b, 160'h5f4c8fa2f113b3637504b42160ddae852daa1d78},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{250, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6e3647dfed9c5ae3cc481528a35f5741e9dc10c1, 160'h569c3937c0a118cb49358a640670916ba346db03},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{252, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h1da6db19788b81fc3ddb980bdefa9a54d33717d0, 160'h018b151eeb8c79bf5be669f12cb784615e098317},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{256, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h3c2c6830a0733d25facdf0048a9d6c3b2921aecf, 160'h0c7e0c333dc82930f5f8a4337b379db7f0a526ee},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{260, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h53a8f7b311fbd2b71cfbc781c50923bf4c423335, 160'h33cf2cf617f565b831d82e93e8fb58de938dbbb5},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{261, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h3332e2dd4080616b964e7bfd569e7b3ca0767b38, 160'h65e0c755d4dcf460fbbd2640d347298f2a29c156},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{269, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h41d8153033a3144823afc2301780de5cc70792fa, 160'h0a9add978d502c71a16a0432451513c7255a4ec4},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{273, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6f10822c847280ca0c687e209d7738db57315dfc, 160'h7ffbab843768815a87be79b2f1edce6be8423480},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{285, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6b7b7ebfcc4acfcb41a8a6a072b745f274382b76, 160'h38a09a2023d79b6242185529aede41eba8f52332},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{287, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h7bf85d33ccb2308d51017419197e53f24a482f6c, 160'h591cbb3ebb4f1bf6571f17b86d07e5f80c6118e9},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{290, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h2ad7961a2515241e9d8675c05aa6fa1488714a38, 160'h17dea0a256ab4e20c9554c5f5b0c491271fb0689},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{296, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b005b80cb0733576bd27520bf7ac44f28e733718, 160'h09738b9aeb21252938e9a5fa885a4bfa3705e084, 88'h01f4c8f927aed44a752255, 88'h01f4c8f927aed44a752254},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=88b(11B), s=88b(11B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00f0a6c8100e5720ab62dc981061abc4add9a1933c, 160'h3673d536905fbe48defe2b2a8637f38f2e1843c4, 32'h7fffffff, 160'h17644e8c2ec89d185d9167f301adcdedae3f5b35},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h711d5c4035baebc8e46bf09434a8aebbb0f678d0, 168'h008f66aea6922e491d02960c4e1baa2c22bcbad408, 32'h7fffffff, 160'h749adb63d26b6d8f49ae9a5725ade8880d9c9b6c},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b3e8857e27393fb609bb7e4d42bb612704d9eef2, 160'h668439313310a849e17faca660f5f5346e11c1a9, 8'h04, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h1b66bc474c8220de08f3db0fdc984b008828ff5d, 168'h00f94509a6596f822f62580acc988bf962ef9e32b8, 8'h04, 8'h03},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h008ac14539432e062ff2b1f6086926bfc87e342e98, 168'h00bdc182b2ec96ac855f1057cd99731a054067a153, 8'h04, 8'h04},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{302, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4a5c77d11ddaa568733d8a6cb79b497e6a644944, 160'h339c2514eda2e275ceffb9a7fc4c8d0470b37638, 8'h04, 8'h05},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h5094345ff85c68fe99627eede704362af196aecf, 160'h53499a272ceb4668c02b4b11e567eae9709f0618, 16'h0100, 160'h1c3870e1c3870e1c387118f7eb1684277916fdbd},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=16b(2B), s=160b(20B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h5e2bb1e908df355fb09ac567021edbc0d0fd7047, 160'h65ee7405ef872af6f2550c123826058ebc8309fb, 56'h2d9b4d347952cd, 160'h1164a61fc3dfa342ba186e32381b34b324117a46},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=56b(7B), s=160b(20B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00de53fcbfc744edfc6be04af83518829b5fa63016, 168'h009fed2940a16623e8f60eec87c32aed905d25feb7, 104'h1033e67e37b32b445580bf4efb, 160'h4cb34cb34cb34cb34cb3e2bdb53bb3e1d213282c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=104b(13B), s=160b(20B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h366bb0c1db172c0da7a94d6b962b2bfb99db430d, 168'h00adb55cacb92dcf86d7e7373db40159c23c6ad8db, 16'h0100, 160'h382efed3dc7e18cf41aec7248f4e56087f9734a0},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=16b(2B), s=160b(20B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0086e01061fc02e52057346370636a5b5cc3710e72, 168'h00ccfb1063a51118d442d5044cb0ecdade51ab7dd3, 104'h062522bbd3ecbe7c39e93e7c24, 160'h382efed3dc7e18cf41aec7248f4e56087f9734a0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=104b(13B), s=160b(20B)
  '{311, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h07970e499d36b850864ce1d6b00d62cb70e2d2e0, 168'h00e30d4b3c346017c766878f93fcbba65cd80a1f59, 160'h55555555555555555555fc42fdb7e4f1437c60c8, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h07970e499d36b850864ce1d6b00d62cb70e2d2e0, 168'h00e30d4b3c346017c766878f93fcbba65cd80a1f59, 160'h55555555555555555555fc42fdb7e4f1437c60c8, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=8b(1B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b1fc10305d2e83868c9e40e8426896297b7f3e00, 168'h0091a1e1f88d1fb0f95380f19c98f55a0854c6b494, 160'h55555555555555555555fc42fdb7e4f1437c60c5, 160'h55555555555555555555fc42fdb7e4f1437c60c5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2b9e690b79e165b04e0df6fc84e58ac94ac63a92, 160'h7a9532b9ee40bff794f9888b1a2e0b8a30f4f550, 32'h7ffffffd, 160'h7ce6e1f81fbdb6ebf382414e62c1c14200249a82},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h409c92512c25d7fdf331487d4bb1ca8312ea27b4, 168'h00db6909d4a0768e609a52064c266e152a36b49b7a, 32'h7ffffffd, 160'h304d26aa02922e73b2c60f12e7f288b0b43f3783},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h39226e3be69faee8861f1fbaf4523da7bd2d1bcd, 168'h00c7a528956daf7f7e5c21288732c69372ca327ecd, 32'h7ffffffd, 160'h2b9afe309194473695a328cfe89a314ee772f616},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h74a34455bc9222dc9f189672e0c72cb3d7bf8491, 160'h605793269a796edfb97deeb50f30477571c76d32, 32'h7ffffffd, 160'h0b63c499d27b74e8894b705f6dcab0b5834c4785},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b1031e0781fecf813633cb3884e930913e65ba5b, 168'h00cc8860779ca7e174df787d66f671a8fa337994cf, 32'h7ffffffd, 160'h3c499d27b74e8894b5a1effb88d50da2d531e626},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00987ff07d407ee7a41a65a7ac6929c13d0a6e4800, 160'h59813e21d5f2fe748f06be7328a9862af2bc7c57, 32'h7ffffffd, 160'h78933a4f6e9d11296b43dff711aa1b45aa63cc4c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h52c0322e296d02806a55800e67b9334ed4005cd1, 168'h00f60f5556e7563b756d8a17cd6977cdde16531660, 32'h7ffffffd, 160'h44a5ad0bd0636d9e12be92d365050cf0ca3e3a94},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50c07170fdea6845c09c3da29cc8ee6700592919, 168'h0099d3cf10ef65514e890c056a08c505ad13dbfe03, 32'h7ffffffd, 160'h15cd7f1848ca239b4ad19467f44d18a773b97b0b},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e2cada2f22ae694fee3a3287ce8dc0691af40c9f, 168'h00f6a592e8c723bec635a76c9c6482d2b60dddb986, 32'h7ffffffd, 160'h5d0e82e246fc758108ac747e6f91ebfc3800d367},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{335, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h009ae2a06f674401b28a799181ad23badd115066d1, 160'h3430009efd1271ea1962d35effebfdf5c94d46d2, 32'h7ffffffd, 160'h44bdeb62114743cb00008678e702d02fe3b75eb7},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4148e9ba110487844c41c6a990ce6029fbacd7da, 168'h00abf5a94d89ac5ad633a85b6879affc41860f2ac5, 32'h7ffffffd, 160'h114743cb00000000000021ccc0e671308267fdb2},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{339, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6f690efb076a7dda2a0f990736ba6cd208144f1b, 168'h00abfccb16e59dd7aecddb51f4e4d2bfc2ae172f0a, 32'h7ffffffd, 160'h67063e7063e7063e7064b08f5189b9de97b88155},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0096d267106dd68444ae300966bac62e18238042d4, 160'h5111e87654afbbad4272a264a6ba5a3320eedc2b, 32'h7ffffffd, 160'h55555555555555555555fc42fdb7e4f118d1b61e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{346, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c1329e5abc05dc8cb22c6c5e900c119fe700880b, 168'h0089643fbd2f156366b3a44316c8bb10e46e305055, 8'h01, 160'h55555555555555555555fc42fdb7e4f1437c60c7},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{348, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c9f7e7bc377bffc4e2a79e4836e61ed5c775dabe, 160'h073a1e62494b22fa27642f51d6f4c5d35d70db5a, 160'h55555555555555555555fc42fdb7e4f1437c60c7, 160'h33333333333333333333975b6507efc3f54aa077},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2102b319abe9060e9d4520b0b6a8ab9641b3b5d3, 160'h2b4067358970714a0f24ae1f351884a7d8588042, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h55555555555555555555fc42fdb7e4f1437c60c7},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a185a284dc8e55e796e084ca5f4ddf5bb8d70a0b, 168'h00d39ec502b4b767c9697963ec98bcd6d613c135e8, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4549f25af5fc3a560c62f91fd555f922df271103, 160'h42890b6465457119a56148c7637a21144cac650b, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h33333333333333333333975b6507efc3f54aa078},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h179d0a5fa8be0b89d8efd25948e8624e3eb1b8a0, 168'h00f614fbdda7c63019c4ad480b01a6f38b7d173138, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h0eb00091546e2d1fc7dcc249da653f08707af318},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00aa5cb12acdf9a8336864190c1dd6df86f98f4c4f, 168'h00b2ffdde9e2b9b558c9bfdf7aa9c7f7ec090c61d2, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h55555555555555555555fc42fdb7e4f1437c60c7},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4f052d5ded4b999f95025401553e1cd6a3f47d6b, 160'h4b4c60ab8e9ab5a0fb004224047396052236b818, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h747c6174595d49f17bb3a36c8b7166421fff8f9f, 160'h5d9784617bdd66817754e964a1c622c40cfdab3c, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h33333333333333333333975b6507efc3f54aa078},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4d0bdafb33dfb43af69e8e130dd901d129ac427a, 160'h1f74bde4f32ad5bb21ae7cae079c9fc583fe196d, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h0eb00091546e2d1fc7dcc249da653f08707af318},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{365, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 168'h00b0046a56f874d30ea2ba7ac1a935fd9d754ee641, 160'h7b9a54d275806819ec30b15618f5625115241f46, 160'h49c9656cd8cbee4456548d63a7fc480791909c42, 160'h6ff78980793ee086a2e66e01a490bdfc03f2d302},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{367, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b0046a56f874d30ea2ba7ac1a935fd9d754ee641, 160'h7b9a54d275806819ec30b15618f5625115241f46, 160'h2dfc21da5c39d441fc6683e54da009f413a0ff87, 160'h647382b3e39a8ac8cbe02f4666d045928a0eb061}  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
};
`endif // WYCHERPROOF_SECP160R1_SHA256_SV
