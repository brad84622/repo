`ifndef WYCHERPROOF_SECP256R1_SHA256_SV
`define WYCHERPROOF_SECP256R1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp256r1_sha256;

localparam int TEST_VECTORS_SECP256R1_SHA256_NUM = 86;

ecdsa_vector_secp256r1_sha256 test_vectors_secp256r1_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 256'h4cd60b855d442f5b3c7b11eb6c4e0ae7525fe710fab9aa7c77a67f79e6fadd76},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 256'hb329f479a2bbd0a5c384ee1493b1f5186a87139cac5df4087c134b49156847db},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{115, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=0b(0B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 256'h00b329f479a2bbd0a5c384ee1493b1f5186a87139cac5df4087c134b49156847},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 256'hb329f47aa2bbd0a4c384ee1493b1f518ada018ef05465583885980861905228a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{143, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 256'h4cd60b865d442f5a3c7b11eb6c4e0ae79578ec6353a20bf783ecb4b6ea97b825},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{230, 1'b1, 256'h70239dd877f7c944c422f44dea4ed1a52f2627416faf2f072fa50c772ed6f807, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h64a1aab5000d0e804f3e2fc02bdee9be8ff312334e2ba16d11547c97711c898e, 256'h6af015971cc30be6d1a206d4e013e0997772a2f91d73286ffd683b9bb2cf4f1b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{231, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h16aea964a2f6506d6f78c81c91fc7e8bded7d397738448de1e19a0ec580bf266, 256'h252cd762130c6667cfe8b7bc47d27d78391e8e80c578d1cd38c3ff033be928e9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{233, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h73b3c90ecd390028058164524dde892703dce3dea0d53fa8093999f07ab8aa43, 256'h2f67b0b8e20636695bb7d8bf0a651c802ed25a395387b5f4188c0c4075c88634},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{235, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h204a9784074b246d8bf8bf04a4ceb1c1f1c9aaab168b1596d17093c5cd21d2cd, 256'h51cce41670636783dc06a759c8847868a406c2506fe17975582fe648d1d88b52},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{242, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3b2cbf046eac45842ecb7984d475831582717bebb6492fd0a485c101e29ff0a8, 256'h4c9b7b47a98b0f82de512bc9313aaf51701099cac5f76e68c8595fc1c1d99258},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{243, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h30c87d35e636f540841f14af54e2f9edd79d0312cfa1ab656c3fb15bfde48dcf, 256'h47c15a5a82d24b75c85a692bd6ecafeb71409ede23efd08e0db9abf6340677ed},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{244, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h38686ff0fda2cef6bc43b58cfe6647b9e2e8176d168dec3c68ff262113760f52, 256'h067ec3b651f422669601662167fa8717e976e2db5e6a4cf7c2ddabb3fde9d67d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{245, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h44a3e23bf314f2b344fc25c7f2de8b6af3e17d27f5ee844b225985ab6e2775cf, 256'h2d48e223205e98041ddc87be532abed584f0411f5729500493c9cc3f4dd15e86},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{246, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ded5b7ec8e90e7bf11f967a3d95110c41b99db3b5aa8d330eb9d638781688e9, 256'h7d5792c53628155e1bfc46fb1a67e3088de049c328ae1f44ec69238a009808f9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{252, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ec9760122db98fd06ea76848d35a6da442d2ceef7559a30cf57c61e92df327e, 256'h7ab271da90859479701fccf86e462ee3393fb6814c27b760c4963625c0a19878},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{253, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h54e76b7683b6650baa6a7fc49b1c51eed9ba9dd463221f7a4f1005a89fe00c59, 256'h2ea076886c773eb937ec1cc8374b7915cfd11b1c1ae1166152f2f7806a31c8fd},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{254, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5291deaf24659ffbbce6e3c26f6021097a74abdbb69be4fb10419c0c496c9466, 256'h65d6fcf336d27cc7cdb982bb4e4ecef5827f84742f29f10abf83469270a03dc3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{259, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5694a6f84b8f875c276afd2ebcfe4d61de9ec90305afb1357b95b3e0da43885e, 256'h0dffad9ffd0b757d8051dec02ebdf70d8ee2dc5c7870c0823b6ccc7c679cbaa4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{261, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h614ea84acf736527dd73602cd4bb4eea1dfebebd5ad8aca52aa0228cf7b99a88, 256'h737cc85f5f2d2f60d1b8183f3ed490e4de14368e96a9482c2a4dd193195c902f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{263, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h499625479e161dacd4db9d9ce64854c98d922cbf212703e9654fae182df9bad2, 256'h42c177cf37b8193a0131108d97819edd9439936028864ac195b64fca76d9d693},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{267, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h352ecb53f8df2c503a45f9846fc28d1d31e6307d3ddbffc1132315cc07f16dad, 256'h1348dfa9c482c558e1d05c5242ca1c39436726ecd28258b1899792887dd0a3c6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{268, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4a40801a7e606ba78a0da9882ab23c7677b8642349ed3d652c5bfa5f2a9558fb, 256'h3a49b64848d682ef7f605f2832f7384bdc24ed2925825bf8ea77dc5981725782},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{276, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h677b2d3a59b18a5ff939b70ea002250889ddcd7b7b9d776854b4943693fb92f7, 256'h6b4ba856ade7677bf30307b21f3ccda35d2f63aee81efd0bab6972cc0795db55},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{278, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h43dfccd0edb9e280d9a58f01164d55c3d711e14b12ac5cf3b64840ead512a0a3, 256'h1dbe33fa8ba84533cd5c4934365b3442ca1174899b78ef9a3199f49584389772},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{279, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5b09ab637bd4caf0f4c7c7e4bca592fea20e9087c259d26a38bb4085f0bbff11, 256'h45b7eb467b6748af618e9d80d6fdcd6aa24964e5a13f885bca8101de08eb0d75},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{282, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7673f8526748446477dbbb0590a45492c5d7d69859d301abbaedb35b2095103a, 256'h3dc70ddf9c6b524d886bed9e6af02e0e4dec0d417a414fed3807ef4422913d7c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{283, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7f085441070ecd2bb21285089ebb1aa6450d1a06c36d3ff39dfd657a796d12b5, 256'h249712012029870a2459d18d47da9aa492a5e6cb4b2d8dafa9e4c5c54a2b9a8b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{289, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4201b4272944201c3294f5baa9a3232b6dd687495fcc19a70a95bc602b4f7c05, 264'h0095c37eba9ee8171c1bb5ac6feaf753bc36f463e3aef16629572c0c0a8fb0800e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h27b4577ca009376f71303fd5dd227dcef5deb773ad5f5a84360644669ca249a5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{290, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a71af64de5126a4a4e02b7922d66ce9415ce88a4c9d25514d91082c8725ac957, 256'h5d47723c8fbe580bb369fec9c2665d8e30a435b9932645482e7c9f11e872296b, 8'h05, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{291, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6627cec4f0731ea23fc2931f90ebe5b7572f597d20df08fc2b31ee8ef16b1572, 256'h6170ed77d8d0a14fc5c9c3c4c9be7f0d3ee18f709bb275eaf2073e258fe694a5, 8'h05, 8'h03},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{292, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5a7c8825e85691cce1f5e7544c54e73f14afc010cb731343262ca7ec5a77f5bf, 264'h00ef6edf62a4497c1bd7b147fb6c3d22af3c39bfce95f30e13a16d3d7b2812f813, 8'h05, 8'h05},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{293, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00cbe0c29132cd738364fedd603152990c048e5e2fff996d883fa6caca7978c737, 256'h70af6a8ce44cb41224b2603606f4c04d188e80bff7cc31ad5189d4ab0d70e8c1, 8'h05, 8'h06},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{302, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008aeb368a7027a4d64abdea37390c0c1d6a26f399e2d9734de1eb3d0e19373874, 256'h05bd13834715e1dbae9b875cf07bd55e1b6691c7f7536aef3b19bf7a4adf576d, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008aeb368a7027a4d64abdea37390c0c1d6a26f399e2d9734de1eb3d0e19373874, 256'h05bd13834715e1dbae9b875cf07bd55e1b6691c7f7536aef3b19bf7a4adf576d, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{304, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b533d4695dd5b8c5e07757e55e6e516f7e2c88fa0239e23f60e8ec07dd70f287, 256'h1b134ee58cc583278456863f33c3a85d881f7d4a39850143e29d4eaf009afe47, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f50d371b91bfb1d7d14e1323523bc3aa8cbf2c57f9e284de628c8b4536787b86, 264'h00f94ad887ac94d527247cd2e7d0c8b1291c553c9730405380b14cbb209f5fa2dd, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h68ec6e298eafe16539156ce57a14b04a7047c221bafc3a582eaeb0d857c4d946, 264'h0097bed1af17850117fdb39b2324f220a5698ed16c426a27335bb385ac8ca6fb30, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d8adc00023a8edc02576e2b63e3e30621a471e2b2320620187bf067a1ac1ff32, 256'h33e2b50ec09807accb36131fff95ed12a09a86b4ea9690aa32861576ba2362e1, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h44a5ad0ad0636d9f12bc9e0a6bdd5e1cbcb012ea7bf091fcec15b0c43202d52e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3623ac973ced0a56fa6d882f03a7d5c7edca02cfc7b2401fab3690dbe75ab785, 264'h008db06908e64b28613da7257e737f39793da8e713ba0643b92e9bb3252be7f8fe, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{313, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d0bc472e0d7c81ebaed3a6ef96c18613bb1fea6f994326fbe80e00dfde67c7e9, 264'h00986c723ea4843d48389b946f64ad56c83ad70ff17ba85335667d1bb9fa619efd, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h03ffcabf2f1b4d2a65190db1680d62bb994e41c5251cd73b3c3dfc5e5bafc035},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a0a44ca947d66a2acb736008b9c08d1ab2ad03776e02640f78495d458dd51c32, 256'h6337fe5cf8c4604b1f1c409dc2d872d4294a4762420df43a30a2392e40426add, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h4dfbc401f971cd304b33dfdb17d0fed0fe4c1a88ae648e0d2847f74977534989},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5eca1ef4c287dddc66b8bccf1b88e8a24c0018962f3c5e7efa83bc1a5ff6033e, 256'h5e79c4cb2c245b8c45abdce8a8e4da758d92a607c32cd407ecaef22f1c934a71, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h788048ed39a5ffa77bfb62fa1fda2257742bf35d128fb3459f2a0c909ee86f91},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5caaa030e7fdf0e4936bc7ab5a96353e0a01e4130c3f8bf22d473e317029a47a, 264'h00deb6adc462f7058f2a20d371e9702254e9b201642005b3ceda926b42b178bef9, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h476d9131fd381bd917d0fed112bc9e0a5924b5ed5b11167edd8b23582b3cb15e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3fd6a1ca7f77fb3b0bbe726c372010068426e11ea6ae78ce17bedae4bba86ced, 256'h03ce5516406bf8cfaab8745eac1cd69018ad6f50b5461872ddfc56e0db3c8ff4, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h357cfd3be4d01d413c5b9ede36cba5452c11ee7fe14879e749ae6a2d897a52d6},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h009cb8e51e27a5ae3b624a60d6dc32734e4989db20e9bca3ede1edf7b086911114, 264'h00b4c104ab3c677e4b36d6556e8ad5f523410a19f2e277aa895fc57322b4427544, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h29798c5c0ee287d4a5e8e6b799fd86b8df5225298e6ffc807cd2f2bc27a0a6d8},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a3e52c156dcaf10502620b7955bc2b40bc78ef3d569e1223c262512d8f49602a, 256'h4a2039f31c1097024ad3cc86e57321de032355463486164cf192944977df147f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h0b70f22c781092452dca1a5711fa3a5a1f72add1bf52c2ff7cae4820b30078dd},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f19b78928720d5bee8e670fb90010fb15c37bf91b58a5157c3f3c059b2655e88, 264'h00cf701ec962fb4a11dcf273f5dc357e58468560c7cfeb942d074abd4329260509, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h16e1e458f021248a5b9434ae23f474b43ee55ba37ea585fef95c90416600f1ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0083a744459ecdfb01a5cf52b27a05bb7337482d242f235d7b4cb89345545c90a8, 264'h00c05d49337b9649813287de9ffe90355fd905df5f3c32945828121f37cc50de6e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h2252d6856831b6cf895e4f0535eeaf0e5e5809753df848fe760ad86219016a97},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h67e6f659cdde869a2f65f094e94e5b4dfad636bbf95192feeed01b0f3deb7460, 264'h00a37e0a51f258b7aeb51dfe592f5cfd5685bbe58712c8d9233c62886437c38ba0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffffaaaaaaaaffffffffffffffffe9a2538f37b28a2c513dee40fecbb71a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0091b9e47c56278662d75c0983b22ca8ea6aa5059b7a2ff7637eb2975e386ad663, 256'h49aa8ff283d0f77c18d6d11dc062165fd13c3c0310679c1408302a16854ecfbd, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h66755a00638cdaec1c732513ca0234ece52545dac11f816e818f725b4f60aaf2},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f3ec2f13caf04d0192b47fb4c5311fb6d4dc6b0a9e802e5327f7ec5ee8e4834d, 264'h00f97e3e468b7d0db867d6ecfe81e2b0f9531df87efdb47c1338ac321fefe5a432, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h55a00c9fcdaebb6032513ca0234ecfffe98ebe492fdf02e48ca48e982beb3669},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00836f33bbc1dc0d3d3abbcef0d91f11e2ac4181076c9af0a22b1e4309d3edb276, 264'h009ab443ff6f901e30c773867582997c2bec2b0cb8120d760236f3a95bbe881f75, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h266666663bbbbbbbe6666666666666665b37902e023fab7c8f055d86e5cc41f4},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008651ce490f1b46d73f3ff475149be29136697334a519d7ddab0725c8d0793224, 264'h00e11c65bd8ca92dc8bc9ae82911f0b52751ce21dd9003ae60900bd825f590cc28, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffff55555555ffffffffffffffffd344a71e6f651458a27bdc81fd976e37},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{337, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6d8e1b12c831a0da8795650ff95f101ed921d9e2f72b15b1cdaca9826b9cfc6d, 264'h00ef6d63e2bc5c089570394a4bc9f892d5e6c7a6a637b20469a58c106ad486bf37, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h3fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192aa},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0ae580bae933b4ef2997cbdbb0922328ca9a410f627a0f7dff24cb4d920e1542, 264'h008911e7f8cc365a8a88eb81421a361ccc2b99e309d8dcd9a98ba83c3949d893e3, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5d8ecd64a4eeba466815ddf3a4de9a8e6abd9c5db0a01eb80343553da648428f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{341, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6adda82b90261b0f319faa0d878665a6b6da497f09c903176222c34acfef72a6, 256'h47e6f50dcc40ad5d9b59f7602bb222fad71a41bf5e1f9df4959a364c62e488d9, 8'h01, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=8b(1B), s=256b(32B)
  '{343, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00dd86d3b5f4a13e8511083b78002081c53ff467f11ebd98a51a633db76665d250, 256'h45d5c8200c89f2fa10d849349226d21d8dfaed6ff8d5cb3e1b7e17474ebc18f7, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{344, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4fea55b32cb32aca0c12c4cd0abfb4e64b0f5a516e578c016591a93f5a0fbcc5, 264'h00d7d3fd10b2be668c547b212f6bb14c88f0fecd38a8a4b2c785ed3be62ce4b280, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{347, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f6417c8a670584e388676949e53da7fc55911ff68318d1bf3061205acb19c48f, 264'h008f2b743df34ad0f72674acb7505929784779cd9ac916c3669ead43026ab6d43f, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{348, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h501421277be45a5eefec6c639930d636032565af420cf3373f557faa7f8a0643, 264'h008673d6cb6076e1cfcdc7dfe7384c8e5cac08d74501f2ae6e89cad195d0aa1371, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0d935bf9ffc115a527735f729ca8a4ca23ee01a4894adf0e3415ac84e808bb34, 256'h3195a3762fea29ed38912bd9ea6c4fde70c3050893a4375850ce61d82eba33c5, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5e59f50708646be8a589355014308e60b668fb670196206c41e748e64e4dca21, 256'h5de37fee5c97bcaf7144d5b459982f52eeeafbdf03aacbafef38e213624a01de, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3d0bc7ed8f09d2cb7ddb46ebc1ed799ab1563a9ab84bf524587a220afe499c12, 264'h00e22dc3b3c103824a4f378d96adb0a408abf19ce7d68aa6244f78cb216fa3f8df, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a6c885ade1a4c566f9bb010d066974abb281797fa701288c721bcbd23663a9b7, 256'h2e424b690957168d193a6096fc77a2b004a9c7d467e007e1f2058458f98af316, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008d3c2c2c3b765ba8289e6ac3812572a25bf75df62d87ab7330c3bdbad9ebfa5c, 256'h4c6845442d66935b238578d43aec54f7caa1621d1af241d4632e0b780c423f5d, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{357, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'h44a5ad0ad0636d9f12bc9e0a6bdd5e1cbcb012ea7bf091fcec15b0c43202d52e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{359, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'h44a5ad0ad0636d9f12bc9e0a6bdd5e1cbcb012ea7bf091fcec15b0c43202d52e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{365, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h0fe774355c04d060f76d79fd7a772e421463489221bf0a33add0be9b1979110b, 256'h500dcba1c69a8fbd43fa4f57f743ce124ca8b91a1f325f3fac6181175df55737},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{367, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h664eb7ee6db84a34df3c86ea31389a5405badd5ca99231ff556d3e75a233e73a, 256'h59f3c752e52eca46137642490a51560ce0badc678754b8f72e51a2901426a1bd},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{370, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h1158a08d291500b4cabed3346d891eee57c176356a2624fb011f8fbbf3466830, 256'h228a8c486a736006e082325b85290c5bc91f378b75d487dda46798c18f285519},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{374, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'h5eb9c8845de68eb13d5befe719f462d77787802baff30ce96a5cba063254af78, 256'h2c026ae9be2e2a5e7ca0ff9bbd92fb6e44972186228ee9a62b87ddbe2ef66fb5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{376, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h766456dce1857c906f9996af729339464d27e9d98edc2d0e3b760297067421f6, 256'h402385ecadae0d8081dccaf5d19037ec4e55376eced699e93646bfbbf19d0b41},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{380, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h6b01332ddb6edfa9a30a1321d5858e1ee3cf97e263e669f8de5e9652e76ff3f7, 256'h5939545fced457309a6a04ace2bd0f70139c8f7d86b02cb1cc58f9e69e96cd5a},  // lens: hash=256b(32B), x=232b(29B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{382, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h31230428405560dcb88fb5a646836aea9b23a23dd973dcbe8014c87b8b20eb07, 256'h0f9344d6e812ce166646747694a41b0aaf97374e19f3c5fb8bd7ae3d9bd0beff},  // lens: hash=256b(32B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{386, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h341c1b9ff3c83dd5e0dfa0bf68bcdf4bb7aa20c625975e5eeee34bb396266b34, 256'h72b69f061b750fd5121b22b11366fad549c634e77765a017902a67099e0a4469}  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
};
`endif // WYCHERPROOF_SECP256R1_SHA256_SV
