`ifndef WYCHERPROOF_SECP224R1_SHA256_SV
`define WYCHERPROOF_SECP224R1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224r1_sha256;

localparam int TEST_VECTORS_SECP224R1_SHA256_NUM = 253;

ecdsa_vector_secp224r1_sha256 test_vectors_secp224r1_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 232'h009e82950ebe102f37ff3645cc7d3c1bab8864e5e03a5011eeba8150bc},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{92, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a040000, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=240b(30B), s=224b(28B)
  '{93, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 240'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad9810000},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=240b(30B)
  '{97, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a040500, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=240b(30B), s=224b(28B)
  '{98, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 240'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad9810500},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=240b(30B)
  '{113, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 0, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=0b(0B), s=224b(28B)
  '{114, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 0},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=0b(0B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h38de5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{118, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h637d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{119, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a84, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{120, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad901},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=216b(27B), s=224b(28B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'hde5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=216b(27B), s=224b(28B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 216'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=216b(27B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 216'h7d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=216b(27B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 232'hff617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=224b(28B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{131, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h013ade5c0624a5677ed7b6450d941fd283098d8a004fc718e2e7e6b441, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{132, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff3ade5c0624a5677ed7b6450d9421a53d481ba984280cc6582f2e5fc7, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'hc521a3f9db5a98812849baf26bdf441fd72b663dc4161062747575fc, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c521a3f9db5a98812849baf26bde5ac2b7e4567bd7f339a7d0d1a039, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hfec521a3f9db5a98812849baf26be02d7cf67275ffb038e71d18194bbf, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{136, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h013ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c521a3f9db5a98812849baf26bdf441fd72b663dc4161062747575fc, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{138, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 232'h01617d6af141efd0c800c9ba3382c2119a390cfa9bed6a409bfe3703be},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 232'hff617d6af141efd0c800c9ba3382c3e454779b1a1fc5afee11457eaf44},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{140, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h9e82950ebe102f37ff3645cc7d3d0508a7abf5a22672e8a95e25267f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{141, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 232'hfe9e82950ebe102f37ff3645cc7d3dee65c6f305641295bf6401c8fc42},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{142, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 232'h01617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{143, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 232'h009e82950ebe102f37ff3645cc7d3d0508a7abf5a22672e8a95e25267f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{158, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{159, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{168, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{169, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{176, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{177, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{178, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{179, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{180, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{184, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{187, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{188, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{189, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{190, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{194, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{195, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{196, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{197, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{198, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{199, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{200, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{201, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{204, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{205, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{206, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{207, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{208, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{209, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{210, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{211, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{214, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{215, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{216, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{217, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{218, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{219, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{220, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{221, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{230, 1'b1, 256'hbacb99f958ccca12280c7b91fb641e03067110ad79ab4268eb8f0786e3f9dbe7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 232'h0096ad91f02a3bc40c118abd416ed5c6203ed7ced0330860d7b88c10ab},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{231, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bcca2365cebdcf7c6cda1ee7b27c7fe79e371537b01869c715eabb1e, 224'h3ae76f9bbfe519d778816dc8fe10635ee7576b6b7916f0c21df320c0},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{232, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h59a9f83289ef6995d5d5592e80ab4f6a81123f69d385d3cfb152faf2, 224'h3a97d5be190d5819241067e2be56375ab84155baab8fc7aeb7f8cb3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{233, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b54bac9be2beaaa09456a3968a1faf27c9d96bd5f6738fec6066d31e, 232'h00d72c22129344a96d52fda60b264cf5e6fae45fd2c1b1b78bcba30070},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{234, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h323dbdecd40910c6fa7a5691846fa7769113d1f2ba64ef0dc97d2ddb, 232'h00ca9e73a4587af042f8ba924bb61829c5e24046f9803eb76ab80ef327},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{235, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a55dccc27d287f15960ed79908a3edb6bb31aff07c8caa0e65fc0785, 224'h559cb51aa5f2b9066610199dd01291a47729a6189a622ae9e7af7621},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{236, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h137ed6105148d6f5b84e87735d57955f81c5914a6e69f55347ade074, 232'h00dfa5d56b1a12567efacb348a133b79d48da7aac78d78ee589c2ec027},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{237, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00856ff63d779163e78fed8c48330b48f08bf953a95266b3857eee91aa, 232'h00f4aa917cd37f556c6df9d0960c2f7daa7ea118e5c30cc40ca1eed418},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{238, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a9d7716f04c5ce247f6b8c608b37db55f68e2ff94a5883863e867708, 224'h61bc093faa6fb25cd240aea4b56fed728f7b3669b4dc84c449d38c5d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{239, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f6d088fd3b9c981ac491c62030643bbd82d4f4588e8517de5884e73d, 224'h773eee477980763b1ea27ae998bda0244cb67b07aa6779a38cd2ba3f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{240, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00eacb55588e446bbf3687089ba8ba3b05cfef7458bb81b4277f90a853, 232'h008039e8944cc3df7f4ce5badc349975d471a81dea14e9bcae3065d410},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{241, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5984af8c89fb9d596a1f28fd3d41e46f7205fe12fa63437ac79e7e81, 224'h33b16b742d45f18f88de2713078384e6150f06b8b99f36ab2ce3dd49},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{242, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3cda62d84711c262f782d5c3a79b567485227b34afb821f5241b1961, 232'h00b615cef399706ff758f072931852b717ec898e9a1e6339d0ee81b8da},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{243, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e1db7304609191ea1ac91183ffb31df51b5b3fdc6b1a1129d85818d6, 224'h441886d003ae80fbe7139e1d02845cd1bd959f0df1468f5836dd6ea5},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{244, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3545dc4a4ef84bbb3a526ff929c91ad234516a9e95455ac8db4012b1, 232'h00af49926f693a7cf11f71e199f382a8d640c0c85e46d94ee26e384344},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{245, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0ccafdeae4582c9de6795b2d09a7fc3848c75904fa960989156cbbb9, 232'h00af1f994da3e7d89cc8aaa44616cb77e3be7a83ccecc965775194e502},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{246, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a3b2145d8c669027532501eea1913abb22a78a827fdd82fe9d6d3757, 232'h009b2f1ae84f5606d68653065f74e9d089886694c739fbe3fd4a1b2b4a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{247, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009aac3a7e3d142344991bf177b4f4dbfa074148ad9e20f27555b547d9, 232'h00f830a3c7fdf251d79d41977d28e6d9a72a36df11b86e17c8dc3acae0},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{248, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4769fba554fd436051c285bdadfa33a443d4f7084dd598ce3b98b8fb, 224'h0c014c87cb14113d75864f74905f75b34f9970ba58b5d0676021826d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{249, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008b91fc5054a75c34a508624b85708b3d25fa74328c68741c3aeb92d9, 224'h155e3e46b1209583135a9fef15abe325b25bd19285ee6b5b4549629f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{250, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a4a2a85fbb8bb26c4d845cfac191f89d65b00d3f1b9450d177f78890, 224'h6605a460e60402685c7a5accd2615e9232e51937bd83dfa3065eabf7},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{251, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a89d333ae34187855cf7fa435ff39be6b7bb39b2d0ce682133ad9646, 224'h483dcc89a3b43be250f5c3f78f78418e7b8341a8bcfb93dfd58e46d8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{252, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2d0f99c71933c82ded544ef4faac9d669e437dea13b57186f4c20a0e, 232'h00d9682b9f3a05d7832947bc45eadbc742d96e7ab1124832ddb7a8c65b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{253, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00840208f7c41b1fbadcc701fb3a1d0f98a3e2a75235e695bfd378f8b4, 224'h44c8daad4efc03e1753803c362b409c3ca6e0f21e538fe3a364c0e53},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{254, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0087cc582cb10602110566fcb10a233aede993fae5fb3f81b0bbff94ca, 232'h00c971c05bd51d9685825b2cfc0a2596c7f80d9f9dc68c28c159aa395a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{255, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h50d73d949b3adcd3e8fa94dafefaf9d263ebc702128d891afac47ea7, 232'h00f8423c378f0190574925142eb5b97c612abfa048fa3ab5375ec795a1},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{256, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d608915dfcd5d3c63ed10d0d9b614f7a866f8858a6e59dc03eb0a8ee, 232'h008e701aa0bab491430f6e4da92244b0bb174957ee6f495bc5d15fabb1},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{257, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c87b0ab842c4769ed94b910bd7719691f9991bc5a347889608f07034, 232'h00d083111048d6e019771fc2669c55156a3d09615a6b2d9cae52ddabee},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{258, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0a1c2c2478e244464226c660edf724db1213f4923eb725d611d976fd, 224'h764e55186a76f734891d05fb57af2727fab8fbea684ca4321d5de540},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{259, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008a2747c5dd9ef5298b8aeabd2fb3a2beb16158fb2cc62be9e51b2152, 232'h00f96251bc048bcad832e6cbc09c9c2e585ab7543dc552eaa5125be0d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{260, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d9eac32a734f3a3e5b5a2905bed8164ef4c6cd24d5c0fc54cc83f3cc, 232'h00a784930d16c3b753bb3ed9151d583c50ff97bc976274bde482fb9644},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{261, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6c40c6b15ae573f77b677cd878cc5e4da8171cf50d79974fde374e00, 232'h00c88c9828037bf7013a1415537ca074d6c8a553bdb4b26b14a7e88d93},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{262, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00dca0aaa0a395393142b323edced09372760350f2ab261ce3339b114d, 224'h0983bf6e510ce7f0a7520f2b7c60cd68a4912b78162c7ac33789e0c6},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{263, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a0526ed47e2607e6bae6dcf3b8f54f4e0638023673a38cad4569c3ba, 224'h61516f55746b379d11cbaa02cef35311d7771a47d1e127cff46dcfd6},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{264, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5c00db60178c8361092bdfb47fc9a47b33363d7e0d76e32520f79657, 232'h00e1baf7ae7d81045793c73173f49d60bdfc8779942795d9d082b3ca11},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{265, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h46f69b6a99717949eee74092a0c1438a290a2cd82fe1e10d8f37e88b, 232'h0099a5f59f09bd980a066233523397846987a8a1bfdde355062d140a4b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{266, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e643d8085a22706fa0e6540f3d5e169ad8cc49b4bfe98e325321c705, 232'h00f95bd423f9cafe0cedfec6fd97871536d71b2ac58dfb2f7ab8952d4b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{267, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e65fb9bcdd791f141ccff2b3cfbf45d84f8c6272021a68dde8c36bc8, 232'h00df6e08c74b5e36b7772658f02515ae0ea813b64df24f3522ea15fb15},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{268, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a476d468221ef55611e8a724c9b4cd79c34f6940d5f665e3335f6231, 232'h00bfddc18e7a008bc206c8e1ca6c878363e4138508e0c3a84a27eabe35},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{269, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1b393477941879271873a8c043a77caadb9957fcdd263a6ac978e4ba, 224'h270060d5f356ebb6d185772baa78b878af6807378e0d5c532da0a4a7},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{270, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b2eda8c969d4b1bdd31867fd1f92d547b406840c257f2f80dfbdc4e3, 232'h00e6297b059ce64ef04de9715a8f686a9f73980865066a94975b7f8117},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{271, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00938189a18a4bff5712ac99c2b8e92c218af3e4d4e3a84b906b0f704e, 224'h7bb3e538f0b70664dad462ab14b0ed416c86ac6e9060fe760dabb715},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{272, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bb7c1d8120d2aa7765b16eeac44282de605fb2a1665657dea4492935, 232'h00e0a8adb3a143883f981ea1323fa6f1d347845be2b8dcc6cd5cc93ee5},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{273, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h74a4c51dd60c7118467be29652060f39af94f8c0eb7f15c64771010c, 224'h6102ec0c9257e607af3f3ff7490b54e78111f422bec11ba01277171f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{274, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h625da18d676f02fae9dbcb3092265909488fb95d662569d7746b9687, 232'h00c4f1ec831e36604d604b630fd0b1999cd09960862294251d85e5873d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{275, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ee0d4a31fd1c4d854d75c14151926899dde1c7332fd4769443d213d, 224'h4b8278b89ba4f8fbd7dcc6affe4c12156f7409909416989685dd5a39},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{276, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdde45fc9ebb3749c9fb2c25bf02e2a217ccc112f8e65499eeffb6a1, 232'h00becd6b88ef2bee872ebc0e2b805a56066e19179fce9f0dc0df3f6378},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{277, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h50186e023a1f5053fcb4d0473039b1b2cdeba569719a4ebabdd675c8, 232'h00f8fb893c1b6b5b827b5f3f4bb5eab75b6212bb56a5a39bb35c127a1c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{278, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d3b454639b0fb3da93b20d55be8609e40902cb4a608f3b9064c0deb7, 232'h00ec7aa9637fd71b543e5243faab4c7a2edc2c48e982c5ac017807f19a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{279, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c202abbd98e03809de842bdef268a1c616a7306da69a87abaf03169c, 224'h7e7e04823af8ed6836fd2ac011e47de8e1bef91ed1da5144893fc259},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{280, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2e4b76638816cce057a4a27a49258dcb5437ae97739f27ebc0973c0b, 232'h00e9f6c0b64e764ad39dd92b576e11c23e5994b02095cb2a4720c8662c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{281, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7e0f48761089aa4c7ecd5a7ac5380836b1e5d381d3400174d15df98b, 224'h0c3df50060e3a6714aa565a33d784e7b16ac87bebfb3c2255cfd832c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{282, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4d6f7408508eb0814dcd48007f0efd9e2b91cdac4030540cc678de19, 224'h1e74f8dc34d13613ef42462fe88981cbe2489be10e4cdae975a1b38e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{283, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00967f2c5d304c7932eaaa1682197945e66cc912b703824776ef16ad7a, 224'h73957001d9037c63d6471c809a2388383ad695137c622cd5f5584414},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{284, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h49260804bb2ceae4b9cee63b02ea60173ec3f4f90167627c0bb39888, 232'h00c9eb022f96db3e90fe0ff617730a629f342e02fb208d6836cbbdc7d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{285, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f3e712597a4b22632c5f8eb9f2845882bb03a139735f80af8826fc56, 224'h62865bd91c0903511a481d607eb6b5fe28f6f6c89295681a3e8d55d8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{286, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0093b4c28f032d00f80e77491edc158359909ee9e30a7327b74219e5e2, 224'h482c19ae35cb28afc9b95ca1ed7ad91c812d5fcceb4beddbf1a16d92, 120'h00e95c1f470fc1ec22d6baa3a3d5c1, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=120b(15B), s=232b(29B)
  '{287, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0093b4c28f032d00f80e77491edc158359909ee9e30a7327b74219e5e2, 224'h482c19ae35cb28afc9b95ca1ed7ad91c812d5fcceb4beddbf1a16d92, 232'h00fffffffffffffffffffffffffffffffefffffffffffffffffffffffe, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{288, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00da927f4ba88b639bf5334221d2f54d8ef9ccc1a1125fad18c7bfb789, 232'h00ac51ae53de6d834a9db3947b8dd4c6ac2b084b85496bfa72d86b6948, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{289, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h20888e1c0f5694c4c0363b36482beb6e1e6649b3d3b26f127febb6fc, 232'h00de00c2f3d8e4a7e8a0bafd417c96d3e81c975946a2f3686aa39d35f1, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{290, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h009545c86f032c5df255a4490bb0b83eca201181792ad74246874db229, 224'h405264c283063327b70f4c2be5ab4d2e9407b866e121d6145d124c04, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 232'h00bf19ab4d3ebf5a1a49d765909308daa88c2b7be3969db552ea30562b},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{291, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h579d53f39d5109bd440e3e3e7efd603740963348ff9c72c03b0fe6b8, 232'h00df02f133ecd60b072a0812adc752708f2be9d8c9ad5953d8c7bf3965, 8'h03, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{292, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d2a14c8106d89f3536faebdafcd4680f65ab4bf2243164ca1464b628, 232'h00acaf2bee52e6231d3c980f52f8e189a41c3e3a05e591195ec864217a, 8'h03, 8'h03},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{293, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e892479153ad13ea5ca45d4c323ebf1fc3cd0cdf787c34306a3f79a4, 224'h326ca9645f2b517608dc1f08b7a84cfc61e6ff68d14f27d2043c7ef5, 8'h03, 8'h04},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{294, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e892479153ad13ea5ca45d4c323ebf1fc3cd0cdf787c34306a3f79a4, 224'h326ca9645f2b517608dc1f08b7a84cfc61e6ff68d14f27d2043c7ef5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a40, 8'h04},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{295, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2b0eac35c0b294f6d435dcaffa8633b0123005465c30080adbcc103a, 232'h00d465a63bfb71d4aee09328697fe1088753646d8369b8dc103217c219, 8'h03, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c6f00c4},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{296, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d156e01e33becede8f4fb4ae9521d751e7f8eb795ca00857db2fd7af, 232'h00d73a450ec60e6a9218a8431870687e0968944f6dc5ffeb30e4693b7c, 16'h0100, 232'h00c993264c993264c993264c99326411d2e55b3214a8d67528812a55ab},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=16b(2B), s=232b(29B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00f293a8a2b4aff0bed95c663b364afe69778d38dd7e7a304f7d3c74e6, 224'h17dfd09e7803c4439a6c075cb579cde652d03f7559ff58846312fa4c, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d4ddf003b298cbaa7d2edc584b28b474a76162ed4b5b0f6222c54317, 232'h00d4e4fe030f178fb4aa4a6d7f61265ecd7ef13c313606b8d341a8b954, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008a5bf0028f1e3eb6841dee7b8f873f68b0c560e592e3182074f51ce8, 232'h009668c32224b65b6849713d35e3acf1786862e65b5a664b47a098caa0, 16'h0100, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=16b(2B), s=232b(29B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b53e569b18e9361567e5713ee69ecbe7949911b0257546a24c3dd137, 232'h00f29a83334cff1c44d8c0c33b6dadb8568c024fa1fbb694cd9e705f5a, 104'h062522bbd3ecbe7c39e93e7c24, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=232b(29B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h77f3ebf52725c809acbb19adf093126a2a3a065ca654c22099c97812, 232'h009f1948d23c5158ec2adff455eb2fedf1075d4ec22d660977424a10f7, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c29bd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{302, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a7f7b99e5cdc6fec8928eff773ccdf3b68b19d43cdb41809e19c60f3, 224'h1736b7a0c12a9c2d706671912915142b3e05c89ef3ad497bd6c34699, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a7f7b99e5cdc6fec8928eff773ccdf3b68b19d43cdb41809e19c60f3, 224'h1736b7a0c12a9c2d706671912915142b3e05c89ef3ad497bd6c34699, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{304, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h009cf00010b4ad86636f6cc70fb58c3b995c0d12e46fc58e24b0d28f69, 224'h21c8a8a320cc450ccb15ebd71617f4ed25db4d3413fbdf157d31dbb6, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00ae9b3636b8547232df438559b5a109e0238a73a76afc25d070ea2742, 224'h7210a69de44ad645b1b03845040f46fce238e92c131a71e4b184c01f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008d57d4fce62757791888c1938076fd766daeb2ec9f1bda8ad5df4809, 232'h00aade924d7ea3ae5abbd0719a7d4865759da654cf76cf7ec031277108, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h10518eb7a926b5f7b65be801ec9b2abf76adce25c6152e452a3512c8, 224'h3f322b9ab57ea8352ad29beb99ef356b713432fcc4aef31f903045d9, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419fe},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008a5dfedc9dd1cb9a439c88b3dd472b2e66173f7866855db6bb6c12fd, 224'h3badfbb8a4c6fd80e66510957927c78a2aa02ecef62816d0356b49c3, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h44a5ad0bd0636d9e12bc9e0a6bdc74bfe082087ae8b61cbd54b8103f},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0083a59fc3df295e84c290b32d0b550a06f99456fc2298e4a68c4f2bff, 224'h1b34f483db30db3a51d8288732c107d8b1a858cd54c3936e1b5c11a4, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h58bada578a205d6e170722c8ed6c7715011fe33d7eba869ed1d448a7, 224'h5be4730c1d2d2ef881e02f028a241b7d7d3b0d0b4a9c0565fcb49977, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaa0f17407b4ad40d3e1b8392e81c29},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{311, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h7fcc799b919fe9789ce01dd9202731cb7d815158bc6cb8468760247c, 224'h0f9d2957e0dd5e4c40124bd5e0dd1be41c038fce2cd1dc814e0af37d, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0093c8c651653430cb4f1675fc86b5e82ca04ff2ab1501674476aac169},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{312, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h3ddd68f69d0bfd47ad19370fa3dc72eb258268c2b5f3768852151674, 232'h00fbe0e155d94d2373a01a5e70f1a105259e7b8b1d2fdf4dba3cf4c780, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h009df50acc33b3625a2d5940dd13dbb97d1f7dd56afff8b7de7545127c},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{313, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h1cb1f564c29ebf60a342b3bc33c8945cb279c6c1a012255c874e1c37, 232'h00b75191ab3b2bb730914ebfa14080410970b71eaf4fe01e2d48be9891, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00dce8c223f235699d1f5d2dcde4809d013390b59129f783239525c08f},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h44e309eb686e7af7f1e2cc17fd56542b38910b3b7908ea54fb038d36, 224'h477e829d4c8332e5b29f344ad27a21c18dab24a31ce7985b63a21304, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h074aae944ee7a7d544a5ad0bd06366f872d2250ba3018a63d2a7f2e6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c728064542cb5142f5eefe638124dcd7a1ad0b3555842a47dd5108e1, 224'h10129dd878ebd47313276cec86f521ea9585cd105b3dc421141993b8, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00aae944ee7a7d544a5ad0bd0636d9455f4e83de0f186f89bca56b3c5c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c46c1ad3d3d0df8e9c0f525c21ce8d81ef9d66297f442d6309966722, 224'h0cfa2253aa31a98d8966b85969bf9c819c019292ef6a53ac1db2a108, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h55d289dcf4faa894b5a17a0c6db3741bbc4ecbe01d01ea33ee7a4e7b},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b7b2e48c1e60e20925f4d9b6be600dd83786a936c9bfab00639c33ca, 232'h00a967cbc65070739a3379da80d54843a18d9c11a29a32234a0b303c12, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h4ee7a7d544a5ad0bd0636d9e12bc561ce04faaf1312bba3a15601ebc},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00f4a3d4598875af7f2741bbd67b1733b6541bc5325b3bcb4d3267c27e, 232'h00c30bf322f58a45c6c2aa2ced55f175d1cbf72a7c5bfc464d74f666c0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h361b9cd74d65e79a5874c501bca4973b20347ec97f6de10072d8b46a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h56d1e5c1d664f6ce2fc1fcb937a7ce231a29486abf36c73f77a2bd11, 224'h6cb282c9d7c6fc05f399c183e880ea362edf043cd28ffac9f94f2141, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c3739ae9acbcf34b0e98a0379492e764068fd92fedbc200e5b168d4},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h30bce8c6b7f1bbba040b8d121d85d55167ac99b2e2cf1cfac8b018b5, 232'h00f1c384c35be0ae309a5cb55aba982343d2125f2d4a559d8c545359cd, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00a252d685e831b6cf095e4f0535edc5b1609d7c5c7e49a301588a1d3e},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e87e538a978cf187908beb27a4a247d496a8421dab1fe79f8744d2b5, 224'h539b9f8fe8bddcf7c97c44c55a4fc22f4d78f6a961447a5b613b5c49, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00ee746111f91ab4ce8fae96e6f23fd9d20a24d2e79eea563478c0f566},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h113a2cc57c8ee7de11bc45e14546c72a29725b9a7218114ac31f0281, 224'h6c765b9a46b0215312a3292f5979c98d37b35883baa156281b1bae8c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h23dd9c3f1a4b478b01fa2c5e997d0482073b32918de44be583dcf74a, 232'h00d661a5ed579a2f09d2ff56d6b80f26568d93a237ca6444b0cadc7951, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00855f5b2dc8e46ec428a593f73219cf65dae793e8346e30cc3701309c},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00bbce4b17d45d24a1c80bc8eca98c359d5e1e458058a00b950643256d, 232'h00fe09e092318e39303dca03688e4ecf300300784312d617e5088c584c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h035f58446c1bdbeaa56660a897ebf965f2d18820c7cd0630f04a4953, 224'h47bdfaea60091f405e09929cb2c0e2f6eed53e0871b7fe0cd5a15d85, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0084a6c7513e5f48c07fffffffffff8713f3cba1293e4f3e95597fe6bd},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00911c0033eac46332691cb7920c4950eed57354761e1081a1ea9f1279, 224'h508ebf7cfd3eab5dabdee1be14ce8296b1fc20acfaac16f7824c6002, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{327, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h62b2abb70bb9c7efdfb57181f433b64751f108130dce180d6992e7d3, 224'h124b3aa8a53e5eedf72aa67e6edcc71f19e36e6ad1d099a59ffd9555, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d8ea27cbe9180fffffffffffffff3a43fa3662a899627950d4eb64bc},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h0f759330e7992752aae6a85f7bb0599784bea53e288ff7ee8d53d5e6, 232'h00defe617362380e92f9a23c4fdcc34e09713aab9cc44119418f6f2fd1, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008f2eda42742ab31f5d4cf666892d1d623efd3b26f7df9aa70296e80d, 224'h3beaf235cfea41fadb98c533a8fdeb5841d69ee65f6e71914711f138, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00bfffffffffffffffffffffffffff3d87bb44c833bb384d0f224ccdde},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2bcf4371b319a691ed0e2e0c4a55a8a9b987dec86b863621e97b9c09, 224'h5b8660a74cc964a6af0311edc6b1cd980f9c7bf3a6c9b7f9132a0b2f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a6f252568f6fbd1ae045e602344359c0c216911723748f9a3e7fadec, 224'h3b76efc75ba030bfe7de2ded686991e6183d40241a05b479693c7015, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{332, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a74c1c3a31c7d493ab2c0af89cf5e688621ca9466d2ba1d8761c3fe8, 224'h2ba0d08f4c9f76856c2b7138c8f1e780b6959992b16ccdfd925f4b3a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0096dafb0d7540b93b5790327082635cd8895e1e799d5d19f92b594056},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h034ea72798257f33f24f64c49438fc43e8f67ddc7170fd127e2c43f2, 232'h0080562acc9b49f2d7fcc89421d2a5db2ea8dd0361fb48d897d4612627, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h3f552f1c2b01651edf5902650fe9ab046f71999ac928edc0087bdb13},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{334, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h034ea72798257f33f24f64c49438fc43e8f67ddc7170fd127e2c43f2, 224'h7fa9d53364b60d2803376bde2d5a24d05722fc9e04b727682b9ed9da, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h3f552f1c2b01651edf5902650fe9ab046f71999ac928edc0087bdb13},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{335, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h3672ba9718e60d00eab4295c819ea366a778dd6fd621fa9665259cb6, 224'h7ae5e847eeaea674beeb636379e968f79265502e414a1d444f04ae79, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h33eeefbfc77229136e56b575144863ed90b4c0f8a9e315816d6de648, 224'h051749dd11480c141fb5a1946313163c0141265b68a26216bcb9936a, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{337, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00bda03b24b62243c61e288b6ea1e99a2886f700944eb1b8f0466cffd6, 224'h1c712a3aaace69331989b707e69e8de39d7cd1aeb65d97ad1800bf7f, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h7abba0cbff134ddcf54d04846f954b882ca9faefdfe818898bfb378b, 224'h792f10b57970ae57bb4fb01c08886848855aeb1984d3d6fcb2b412df, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{339, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00f68d99e28653b9ba3e7cedb3b78165f5a54fbe90d4b9f88497977e16, 224'h234da3eaa0178a51b5b0c208ef0818df6f6578793c1af1787026b8da, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{340, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h065d9ef133ce81c2d6b66e928360f9527f8f36b5badd35b5f1093427, 224'h2004852755f77440a0b08b9f165489c0696e8b4981d6d04a285b0fd1, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d6cea09472ede574ce1e0546c9acd0e1cd8cba9b121df29e89d5092e, 232'h0083904ebfb902ea61c987dc0508e0c9a7e563e2609feaf79140ab91d6, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{342, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c520b18003b356094147ee2f9df1178572bed837bd89443b25ebceb8, 224'h0e2e93a998fbbabe82192ea4c85651cf09a95ab0dc2e3d975ee7be98, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{343, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h009dd0b99bb7a830bcc7d55abac42912d525b063c50cf377ca5771a26c, 232'h00a141fccf0793c2ba2469a946c2d4ed26344052c63a6d7e7797ce96c3, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{344, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h3dab9f1b19e715d174a7360920375d569a181f055e66f01391871b6f, 224'h47a6d87c23a5b6a1e3d0a9721302cc02cce35f35dea08e22619be521, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{345, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h56dde1ba58ea31053b2535c66623344c24c72d214af5be6982e89100, 232'h00e771084806143e86f2b31bdaf62280f5b311d0d2bdbb385b20fc6c87, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{346, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0094efe1387fc0447d7dbcb53739a0e4e0ddec181d382caea645b1a612, 224'h4414a6b1c78908d0fa206f8f2de950ad4a14d1ce94d9cddbe32e4601, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{347, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h6286803b952976ee1897013695d3ef2cbb6f977142a042b236572577, 224'h722a6ce9ad3e3fd28e451833496c63b8ab70538877215f204942bf59, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{348, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 232'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419fe, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{349, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h44a5ad0bd0636d9e12bc9e0a6bdc74bfe082087ae8b61cbd54b8103f, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{350, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 232'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419fe, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{351, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h44a5ad0bd0636d9e12bc9e0a6bdc74bfe082087ae8b61cbd54b8103f, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{352, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h0364e7d96832614a80216e730c353534d4bffd2c26649c0b4b0e2628, 232'h008f40064b412fe38c5ba9cf664e6172ed48e6e79f0fe5e31a54985dfc},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{353, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00f4b68df62b9238363ccc1bbee00deb3fb2693f7894178e14eeac596a, 224'h7f51c9451adacd2bcbc721f7df0643d7cd18a6b52064b507e1912f23},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00b2970cdec29c70294a18bbc49985efa33acc0af509c326a3977a35e8, 224'h0cea3ed8ebaaf6ee6aef6049a23cbc39f61fcf8fc6be4bab13385579},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{355, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h7e7b0eb7da8c68a7072b11404ee95a5c407fbfe3d69646802e28ae77, 232'h00d409a2f6bbaae59bb60fc0a092b12fa4e67dc8d088cf19a833322fd6},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{356, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h519bf185ff4635271961fa491be257231deeea9c53a6ede3b4a89ed1, 224'h486bdad484a6a3134e1471cf56a9df0fac50f773b3e37d6f327617d7},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{357, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h09fd644898b7cb5d018b52234e7b4ef2b54789afd0ce9c434e9e5515, 232'h00f19309532164ea2053cae55df7bdcbab536c83ea7bfe6fe10d60c1ab},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{358, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h00ec919d4e283ccf1f71a9e3c0f781a36758d3f38b1b78a87a74288e80, 224'h4c4663044a73c79bd88f0dc245ab1a32f89f06f40a704b31e9fabc51},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{359, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00c51760478447217597ecc6f4001bd45088d53c90f53103608bf88aea, 232'h00a201253aa903f9781e8992101d7171d2dd3a5d48c44d8e1d544cd6d7},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{360, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h76be0112674ec29128823e1af7512e6143872fef30a64e2f1799bd56, 224'h187e503e1a48c27b549fe0a4ce5e581e242c8663fc9efb02d6f2b193},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{361, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h36245ef126b5b51e459f84eaaad5a495061f0471dc8c23f1c5f16282, 224'h39e31d72a06ba8e14fcf95778e07bc16a2628e39449da8857d506edc},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{362, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h258682975df8bca7f203f771ebeb478ef637360c860fc386cfb21745, 224'h7663e70188047e41469a2a35c8c330dd900f2340ba82aafd22962a96},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{363, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h0085c98614f36c0d66f8d87834cae978611b7b4eebf59a46bea1b89ae9, 232'h00d1a18e378dda840e06b60f6279bf0a2231d9fa2d8d2c31e88bc1bdd7},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{364, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00ca7b7432ba41ff2112e1116fffde89bbd68f5ce67fe5513d16c8e6f7, 232'h00e421b7599e0180798acc2006451603cda2db1d582741116e6033ce5f},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{365, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h19397fe5d3ecabf80fc624c1bf379564387517c185087dc97d605069, 224'h33b5773e9aaf6c34cb612cfc81efd3bf9c22224e8c4fa1bfccf5c501},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{366, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h70f24f5c164164bfbb8459aa12a981aa312dbcf00204326ebaaabdc8, 232'h00f5cebee8caedae8662c43501665084b45d2f494fb70d603043543dc4},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{367, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h0bf2d86ecaa8b56aca5e8f8ebcb45081d078a14555b75f5be8e9b132, 232'h009a55b3ce4734849966b5034ccd9b19f76407ee0241c3f58e7b8fc89a},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{368, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00bfc5dc4434cd09369610687d38d2d418b63fd475dea246a456b25a3a, 232'h00b171dfa6cf722f20816370a868785da842b37bac31d7b78e6751fc50},  // lens: hash=256b(32B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{369, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h008fdbe8da646c5642d767c7dbeb3872b1edab6e37365805f0e94ce0a9, 232'h00bcf35ab81222883dd3526cb0cf93138f4687cd0b10c2b0a126385161},  // lens: hash=256b(32B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{370, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00e23a11275848fd4f8b6f4ac4fc305eae981d3b7dc453e5a980c46422, 224'h1a875693f24a03ea1614c4c3bbd0dd7221429f22b337ea7d98348ca4},  // lens: hash=256b(32B), x=224b(28B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{371, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h76645164ff9af3a1a9205fda2eef326d2bffc795dcc4829547fe01dd, 232'h00b65bba503719314b27734dd06b1395d540af8396029b78b84e0149eb},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{372, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h32fa0ca7e07f1f86ac350734994e1f31b6da9c82f93dced2b983c29c, 224'h7b7891282206a45711bdfcb2a102b5d289df84ff5778548603574004},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{373, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h2d5492478ca64e5111dfd8521867b6477b7e78227849ad090b855694, 232'h00a532f5a2fa3594af81cd5928b81b4057da717be5fb42a3a86c68190d},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{374, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h191eee5daf55cd499e8539cb2cff797cfec5d566d2027bf9f8d64693, 232'h00dadfeae8131f64d96b94fd340197caa2bc04818554812feef3343070},  // lens: hash=256b(32B), x=200b(25B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{375, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00e0e2c08180b8a207ee9105a7d379fa112368e8370fa09dfde4a45c45, 232'h00c717bc0860e016e7ce48f8fe6a299b36906a6055adad93b416ce8838},  // lens: hash=256b(32B), x=200b(25B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{376, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h1b919ef93532292743bb2e1b7b4894fd847c6e5de52a08e1b0f2dcfb, 232'h00c2d30d6b7594d8dbd261491ae1d58779505b075b64e5564dc97a418b},  // lens: hash=256b(32B), x=200b(25B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{377, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00e75db49ed33ff2885ea6100cc95b8fe1b9242ea4248db07bcac2e020, 224'h796c866142ae8eb75bb0499c668c6fe45497692fbcc66b37c2e4624f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{378, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h1f81cd924362ec825890307b9b3936e0d8f728a7c84bdb43c5cf0433, 224'h39d3e46a03040ad41ac026b18e0629f6145e3dc8d1e6bbe200c8482b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{379, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h00fda613aa67ca42673ad4309f3f0f05b2569f3dee63f4aa9cc54cf3, 224'h1e5a64b68a37e5b201c918303dc7a40439aaeacf019c5892a8f6d0ce},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{380, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00b932b3f7e6467e1ec7a561f31160248c7f224550a8508788634b53ce, 232'h00a0c5312acf9e801aff6d6fc98550cfa712bbf65937165a36f2c32dc9},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{381, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00e509593fb09245ee8226ce72786b0cc352be555a7486be628f4fd00c, 224'h0b7abde0061b1e07bf13319150a4ff6a464abab636ab4e297b0d7633},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{382, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h6e54f941204d4639b863c98a65b7bee318d51ab1900a8f345eac6f07, 224'h0da5054829214ecde5e10579b36a2fe6426c24b064ed77c38590f25c},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{383, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h0085ea4ab3ffdc992330c0ca8152faf991386bce82877dbb239ba654f6, 224'h0806c6baf0ebea4c1aaa190e7d4325d46d1f7789d550632b70b5fc9b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{384, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h44d53debb646b73485402eab2d099081b97b1243c025b624f0dd67ea, 232'h00e5de789a7d4b77eac6d7bba41658e6e4dc347dabed2f9680c04a6f55},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{385, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h1526eb2f657ebea9af4ca184b975c02372c88e24e835f3f5774c0e12, 224'h1f1ecce38ee52372cb201907794de17b6d6c1afa13c316c51cb07bc7}  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224R1_SHA256_SV
