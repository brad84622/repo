`ifndef WYCHERPROOF_SECP224R1_SHA3256_SV
`define WYCHERPROOF_SECP224R1_SHA3256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224r1_sha3256;

localparam int TEST_VECTORS_SECP224R1_SHA3256_NUM = 72;

ecdsa_vector_secp224r1_sha3256 test_vectors_secp224r1_sha3256 [] = '{
  '{144, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{230, 1'b1, 256'hb2d2232f6d22c49f89c3c3a8a99484abbe828ffe8430eff4b891ec16ea512813, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 224'h7eb5cea4bda67eb17c42fd9e4ef8fc07a386c4d38b8e3fd7ac14e601},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{233, 1'b1, 256'h80e10000000005f3acf7efe73a0182b5f719824bfa118c4925a1e8e0f194add8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h44bf0e8ef31adcf935bfdbdbffb848160ef5d5f97973303503ae43c6, 224'h58194109101107d061575d48aefb8791da1aeca9214fcc4bf9b60dec},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{236, 1'b1, 256'h8b9d7d14000000009051340f34c75a0e78f4a191b3f908bfdaa334f32eb47b51, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h21dd71ac10881ea88296395ab8efbe822c081b5a6d448e6e5d6de917, 224'h3b906e2910ac307a545c7c5e5a4155631be6ded9da8719f4590b5df2},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{237, 1'b1, 256'h432701b4c5000000004e77e86a34ff07f3069a9b547da784a05d7d5d950984c6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3c8dd1c1da01ca7793890cecf967aef7b3199be89973f40f132f47cc, 224'h7030a2afbf16e0200c9b5d9104009881b5667f5c991c3150d5ec0923},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{238, 1'b1, 256'hee4ea2312d5300000000f10e2378adc2459d7728a0eb1c3fa70bf25ffdfc2d9f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1bb538ffd49b566203b3390186d41052e2158bd8cabce482e2bd9cfd, 224'h2621fe8a3ebd93982e7ad1f876e354a56809f8cdaf7289c247a93509},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{239, 1'b1, 256'hb519e0108d975a00000000885c7dca69fda64d70ab959d0a99034d75dd180ce7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0b6b5578395738451e59bc461bfc558b0ffadc75045c4298b00f9539, 216'h3147e9cdce81809e25b10531c59ae3f225c7a7681ff5135cf317bd},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=216b(27B)
  '{242, 1'b1, 256'h88c1ae896d5b1ee1e1280000000051e2c22d970dc99dcebfd57a35be0f5195bb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3a9c3646b7af34c502284ef0070287672dd2b59e2e60f7272d50095c, 224'h561225addbaab4b7bceba248b06dd462779bf1ee3198c2ea417ea42c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{244, 1'b1, 256'haf52ca1d210a9ea8ae35e8fc00000000cec8a7eb3b52686105536d8fc3757f7f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2ffec2697a93f0c4c5a48bec8b15dad327b1b70017e6925fa76b683b, 224'h205dbac588cae4f0ed3b8c7b4101399ce183d38211ed22306d0cda12},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{248, 1'b1, 256'h8b15a9990c7fe432804ea9a57b1c8db8000000000033521f6cd85d48845871b4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h33efa91052f2a89dafd2b06cfa28b0c8243e3cac8246c1aea3cf4e60, 224'h41f964715dd55418a5746f91ecff15b7c6163fb94c18979cf693c21d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{253, 1'b1, 256'h01ca3636d480cdce6ee63cbe3665c7bd88995f000000003f5d61628138af2b7a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0fd7a377de13b55ed9e39abed7153ab72b3864ae00089be6cb39c5ae, 224'h01999722036ba44e9e00574b3de46a7c2af46974f3ce38181cebace1},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{254, 1'b1, 256'he64458ff971279b567c8eb016ac86c39f963cbaa0000000056fbecb71ef3fd7b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h179ff07fe7b684e7231efcb22216709b6c5b64f3e2ab2b6962b7d0e2, 224'h3077af624bfa19a3df87362e3a41ea0e7f904b32c06851cee0f5b6a1},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{255, 1'b1, 256'hb15bafa66eaa8c73cedfc9568ac5a41a5b0a45e38e00000000f88ffd117bf4eb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5d6817bbbcfa633f934456ab5946744128bd0eb7c5bbe6db16e9594d, 224'h73c234f3f23187b318b984d099838ef57873ba6de48bd9fadcd2effe},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{258, 1'b1, 256'h1d29293e1f2113a0eec5780d25200ee18779ad86ca0431390000000088a9c6e0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h10a8cc92e550c816999c0a9bde2b345a2a75c6f66861f060ff2a3742, 224'h6ef54556c7883fc45e8b00638ff76c1f3eeafa895e4f2dce990249fc},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{260, 1'b1, 256'haa2ef39293ec474361e7562735439b835b55d17b130df2421eb200000000fc40, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2c3d2fef2d23ea431f36dd3258127326f83aba9989754fd733931bb0, 224'h64de0f37c334eb07f57e5dcf925a7806f90f1af34c2544cf3d4d9f65},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{263, 1'b1, 256'hfffffffffbda4755bba6de00c2701a0c6fd32c7e4aa1d876140f979cc80f34c6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h254485afee6912f38bffae771553aaf734c779b769e792b2623ab056, 224'h6e599ea2fe87d2228992cea340b14d8872ad3cb2abf35a1f453c7c24},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{266, 1'b1, 256'hd0fab1ffffffffbf5c5a0dc94820af6ed2c80b5411be656e273b963141464e36, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5224c582ac8f7101bf6fe14a9617ca0a9878dbbe026ae230d1e63d0f, 224'h61f0e486a1b7cce228874e7ccb6dc8dc95434afe6dbb7494b9f0e1c9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{268, 1'b1, 256'h4d77a2c899ffffffffb8c2d8566f592706ca04276262ff7cfdba0b2ad6e2a6c4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h74d5a5f801ab103a8de9cefe365753e5e4e24aae88b18ead08f9e7e1, 224'h22195ff2b1dff4f8ef7382a52f177a766a8f839b65b77076850c5edd},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{274, 1'b1, 256'h6162159e82cf80a70b34f2ffffffff193b3c777305a8fc809337cb13014edc7a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h27a2c5db14c60f71c3f08196356ea7094db6559a4c5c7ab097aad799, 224'h755741a777ad419b5c1853bc6f8da89c282a67f71cd1fc3abfe6ef1c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{275, 1'b1, 256'hb35876d301bf4040fac24355ffffffff7fd82e02fe5885a42240d05fff5fc61b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b5c4a2123721cf74e151a3f3d97880d198cd7850a490b3736ed28a4, 224'h4b0107b4c7f32a46315160b39f95d2bec469981960eeaf99f30e8d8b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{276, 1'b1, 256'hc5ae766a399aa8c082a59a4f62ffffffffab6578abad5454b86f0be4e36bedc8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h219a8f9d6701d7b51d82b293d2f0ce4847e13abe9dfe8de426164040, 224'h33623e698063becd8f28445ddb16caedfbe093a2c1d89925c28a12f9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{283, 1'b1, 256'h07fc58409c7cb5c7169a63d09e4de5120132b8ffffffff1f95f5e389535720ac, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h38fa40a57e4a04024c899051cc8080c5261dde66ea59fe532e852013, 224'h3e99d123e596e993d677683bd25889549155edae098e59a29fe7d9cf},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{284, 1'b1, 256'h383dfba6e0aa10f820e15e27374c2eb6996baf43ffffffff66a94ff532236f85, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7f62a985c5bbde0e11e0250a97d73fa38011bb83b6fa2d9836bf5c45, 224'h3bd850832cc305e6b7d9566d36951ac4794b2d08ff712b18b0af6594},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{287, 1'b1, 256'hb291bf1a8c66adc9def9a0a96da478aa1d09e06797adcdffffffff8fb0460842, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h075ceeeaa2ffbe5dc173d84df71145a056500a90f8fb902a24c0d363, 224'h688cefcf26f584f8d598da2b960a512b6b65a425ed536a4bd570cf83},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{291, 1'b1, 256'h1f52ed3bbbeeaa23026b261a17bc00058f2e37cba29772831b7ed9ffffffff02, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2ce15f3bc4f827e2cd5f59b7980f694e91c4b6a7b77c616f17121136, 224'h3f71766ac9e52b98f58a6895112e43b75925183a29a73bd835f95593},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{297, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h1977aac0b91c2b65f580a5f33d8045a3a56e3a3ab48d8613f3ac0844, 232'h00c315f37b48cb771635e16afbca84948b9e4e35690a0990bddc6cab9a, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{299, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h6731bd2f7969febf93fa2382bd4fdc93ddeede8f2deac4c3abf1ce7a, 224'h19516b15727d111c786b39ba11026d25a220b4fe52c5f56fd4ca5dec, 8'h03, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4aa4667eacd6788f17ebde59e78dde177b2b378945ba487d325567d8, 224'h5d887d32e8cf6d5182433d8f81c945b4356d3ebc0e970dd0a9035387, 8'h03, 8'h03},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h0322435ef8557da9306c645a0b614c6f6ce98d859697784cf74f2f23, 232'h00a8cd9e243e9088170133bd81eb6cd28571fcf207509819f443e5bbb5, 8'h03, 8'h04},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{305, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b00ff7e1925b9717903a05d40ce9860ed12ebed8c686e05a9205a976, 224'h110ee94a9a3267ab1565c66cdd5ed2844ccc5c6a7e78e4821b954f98, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{306, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b4f18d031097f179effad146f5fa7e8574e6493dc4133a7e6bff6763, 232'h00b11ad9abcde8a93b78b6bc1f71d96168712263f6fdeb1da9b1193912, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{310, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h009c88d34bcdc70a09bd9cb4aab4e40fa900472d635c4ebd2366e5d4b9, 232'h00ecc54c3d44714953766bbb1257a3580a2aa85170e418969ba3a66841, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{311, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h009c88d34bcdc70a09bd9cb4aab4e40fa900472d635c4ebd2366e5d4b9, 232'h00ecc54c3d44714953766bbb1257a3580a2aa85170e418969ba3a66841, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{312, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00a3ce180bd65ffc76d5502ae806a6b434d7e69b39b1940e44c83604cb, 224'h4150ca512dddf3363897dd8d23f76564412188cc9be77c170dcef4e7, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{313, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h7a1183e83dd8e38b2aef19c9e604a205ecf50abc9ad1b2bf3a062ba9, 224'h35d0ec70d1c66ba124872a47d044b8bb7b6a405b9a9bcce636f9e788, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{314, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h6fbbbfa60d49b603fbc7f6f6c922df0364c03f089af3a288ce4337d5, 224'h28c46eb6f43e9c4f2664ff72d587cd706c620cd718bceb1197482ed9, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00d50a93a475ab04521ca4bc4dcd06872e85fc587a7c56e68a6e94846a, 224'h4511f0bd21af19dff4def09b04bcb20e21ad21e0f8c4a49f21856aa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf7},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{317, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4a8ead5e32234b2a78171bbe3215f1b721f9ae113c7e9711bd44cb28, 224'h15580cc1e9f22a432e8070f700b949ea55cfcd9323589fe1edb06053, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{322, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00e0af4ad4f06a41c72d502d6934c8c3f4b34f062d1cf723b3712c9af3, 224'h4a3d09ffd3506e11669609ea8fe8ee54b30188bc0ad136cdcf73038c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h17688246313d0b42a8ce483b42fb1f0a6217394611f2b177ada94b47},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{324, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00e14fb7fc849de20d33c6c5e6b358f5ba702eb2b9121def8d3deddbdf, 224'h58153c8e0ef0b78993f4d17405c1fe2b20880d40b229f7de51a4d6b3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h1048c627a1685519c907685f668c11b76a11dc9e381d35c5efc14b87},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{325, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00f83a254c07c29022454c43be9bd5e99c630ff7d83206713a1fbfa0fa, 224'h017a0adb068fb28a9418328eac1bc19c6c92c3f1666a773250571a19, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h313d0b42a8ce483b42fb3461047c69e7886089d9f0c0fc2c4d917952},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h23ac1ccb807f76fa99207af67f662fb1ee10f1d5fddb715eafa8ad3d, 232'h00b18eceeb7432c70250f8e92fa990baab18296547fb7901acdd8faf59, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h1c22615f35d488bad614c3cc5578205bd25c0d73ed985e1214d094e1},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{327, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h119d9f0c5f5f6206df598622ec7afc756a0c1c1b3d1133528a7a06cd, 224'h0df17a9164719714488b9ba8021885d4eaa83e8842b11af368d06304, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3844c2be6ba91175ac298798aaf040b7a4b81ae7db30bc2429a129c2},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{328, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h008888ae9b1ab8d57b18468a2c16f8c971a70711c6361a9afe14be4e33, 232'h00af32311a18ef6b965c8f6e252051794a3467de9f58c06a8545b743dc, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h5467241da17d9a30823e4b65006861137714285bc8c91a363e71bea3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{330, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00bae5f11eb77e354a0d0e33c4ce24839d726e1700e514ccbdede23145, 224'h4ffd009fbeea9c7307938f8adfed84de3600920286281d267c88609a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{332, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h39b30cf6827e95c4bb1cf5a201e3611ea87660c671fcfe4837a55ba8, 232'h00bf990d7e7756ab4c0f08f0d674980caa2e559c93c84f7042fbf0ace0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{334, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h69211fb68e0ce40b590bdfb262753d3817a9777cbcc18292f63d9446, 224'h7fc0dcf4d6a02a0daf952f1bdc99ecb4bcefde8d7eb22ae14be44b5f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{336, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h1a51969a30f966894ed0e1b763da7cdd2a258a9a9d6efb019419c152, 232'h00fd8982295489e97f2d8d6ebe0409d759a5ca25cf9627f20e39f1e651, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{338, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eec9dbb6fe5ed5c8e4f8309cd81d506005efd52dca73e8874957db2c, 232'h00840f6693e77f92088c6e411075ff15817ca0f6e669a295d01d2442bd, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{339, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00a4b5e9304fb04bc6257fed45083fc7f50aacffb962d42b3b3a6c6177, 224'h58aa38fe0aa034025e4b7ed045eea3edad0a5ece26bfa7441239f521, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{343, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ebc69137db89c0189696ee75ff03706b0d939639bb64e220d70ecee6, 224'h23a446d65b083da18cb14cb6a9e57f007558386065726ea34feab573, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{344, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ff8f64c0c0f7f0e81d205b67a1c3bccf0c3dcf3bfdfdc80a61471e80, 232'h00a0cbbf29ebedf5381016937ad91335c5801bbe6fd4a1ee6199295601, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{346, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h3e4fa16464ba762f06e7cec2fcbf66269ff742c10a53361217f2053e, 224'h706b308fa36b5de586523d32244eea63a4d86f215930eae2bf99808e, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{348, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h235c610afcdc0a22f84d753b1f7b9cee388f8f5d68127046500b4f1a, 224'h605e49168429c44e190d3612f355bd7e63978fb6c9a61dcd53b13821, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{349, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h009f77906d353c1b862ec4794687c69fa506405c4d0b57f4ef8491dba7, 232'h00ce9e810af65edf1ae583e6f9d6f2ddbc01365e1e744f2987af5527e0, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{356, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{358, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{360, 1'b1, 256'ha7ffc6f8bf1ed76651c14756a061d662f580ff4de43b49fa82d80a4b80f8434a, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h2a8e4fc8c813be0459fe6fd5a449fcd27118121180f37f96857498fb, 224'h487fabaabee79f667da6505c5c171d299732d37784fd73775dfd3db3},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{362, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h295e399cbf4904e22850240598e009d6b40d6391e370aba5a04042d9, 224'h2a0c5841560271a38c7b7c3bb064990e204bae693e2171a246942d40},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{366, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h3e4f9883f7acaadf2a076234fa99fd25a5d8369fb7766aa5b2eb3fd2, 224'h42cb3e2eb9f5431fca4a7ec83637aca92fbebe8afa4ab4bced1088b9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{372, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h4b9b6fefe18c73272ee66ab96fe340b3835b1f63f903b1ac76ba3457, 224'h0c580a65c53b48d1180f0985fe0f9d5f57cf7eb5e572b9714411aa98},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{385, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h3a224d4baaa5d5c332a3d62043b1aaf66b029880010c839c5c033aa3, 224'h2de87b37b0305cf6112e0ac94200118ff493c0a379f4beb0b6602e02},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{388, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h5c7c63a63a69787bfc469ab70a6856f7f322447f9ce74573d0f94d2d, 224'h3e80ff0a9fbd8c11a08d7dc02237e435838de2d2b51eec1156e667d1},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{391, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h1023fa4d5dcedab53a8fdfe2a8f8da941be08c63146e4ba2ed87bd4d, 224'h367a88e393fd1ee4ec925f7f920d4c3fe3ba48edbd253261ec706c5e}  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224R1_SHA3256_SV
