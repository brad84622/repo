`ifndef WYCHERPROOF_SECP256R1_SHA256_P1363_SV
`define WYCHERPROOF_SECP256R1_SHA256_P1363_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp256r1_sha256_p1363;

localparam int TEST_VECTORS_SECP256R1_SHA256_P1363_NUM = 214;

ecdsa_vector_secp256r1_sha256_p1363 test_vectors_secp256r1_sha256_p1363 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 256'h4cd60b855d442f5b3c7b11eb6c4e0ae7525fe710fab9aa7c77a67f79e6fadd76},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{3, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hd45c5740946b2a147f59262ee6f5bc90bd01ed280528b62b3aed5fc93f06f739, 256'hb329f479a2bbd0a5c384ee1493b1f5186a87139cac5df4087c134b49156847db},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{5, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hd45c5741946b2a137f59262ee6f5bc91001af27a5e1117a64733950642a3d1e8, 256'hb329f479a2bbd0a5c384ee1493b1f5186a87139cac5df4087c134b49156847db},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{8, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ba3a8be6b94d5ec80a6d9d1190a436effe50d85a1eee859b8cc6af9bd5c2e18, 256'h4cd60b865d442f5a3c7b11eb6c4e0ae79578ec6353a20bf783ecb4b6ea97b825},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{9, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{10, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{11, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{12, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{13, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{14, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{15, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{16, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{17, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{18, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{19, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{20, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{21, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{22, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{23, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{24, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{25, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{26, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{27, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{28, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{29, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{30, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{31, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{32, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{33, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{34, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{35, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{36, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{37, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{38, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{39, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{40, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{41, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{42, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{43, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{44, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{45, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{46, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{47, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{48, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{49, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{50, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{51, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{52, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{53, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{54, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{55, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{56, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{57, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{58, 1'b1, 256'h70239dd877f7c944c422f44dea4ed1a52f2627416faf2f072fa50c772ed6f807, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h64a1aab5000d0e804f3e2fc02bdee9be8ff312334e2ba16d11547c97711c898e, 256'h6af015971cc30be6d1a206d4e013e0997772a2f91d73286ffd683b9bb2cf4f1b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{59, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h16aea964a2f6506d6f78c81c91fc7e8bded7d397738448de1e19a0ec580bf266, 256'h252cd762130c6667cfe8b7bc47d27d78391e8e80c578d1cd38c3ff033be928e9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{60, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h9cc98be2347d469bf476dfc26b9b733df2d26d6ef524af917c665baccb23c882, 256'h093496459effe2d8d70727b82462f61d0ec1b7847929d10ea631dacb16b56c32},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{61, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h73b3c90ecd390028058164524dde892703dce3dea0d53fa8093999f07ab8aa43, 256'h2f67b0b8e20636695bb7d8bf0a651c802ed25a395387b5f4188c0c4075c88634},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{62, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hbfab3098252847b328fadf2f89b95c851a7f0eb390763378f37e90119d5ba3dd, 256'hbdd64e234e832b1067c2d058ccb44d978195ccebb65c2aaf1e2da9b8b4987e3b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{63, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h204a9784074b246d8bf8bf04a4ceb1c1f1c9aaab168b1596d17093c5cd21d2cd, 256'h51cce41670636783dc06a759c8847868a406c2506fe17975582fe648d1d88b52},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{64, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hed66dc34f551ac82f63d4aa4f81fe2cb0031a91d1314f835027bca0f1ceeaa03, 256'h99ca123aa09b13cd194a422e18d5fda167623c3f6e5d4d6abb8953d67c0c48c7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{65, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h060b700bef665c68899d44f2356a578d126b062023ccc3c056bf0f60a237012b, 256'h8d186c027832965f4fcc78a3366ca95dedbb410cbef3f26d6be5d581c11d3610},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{66, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h9f6adfe8d5eb5b2c24d7aa7934b6cf29c93ea76cd313c9132bb0c8e38c96831d, 256'hb26a9c9e40e55ee0890c944cf271756c906a33e66b5bd15e051593883b5e9902},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{67, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'ha1af03ca91677b673ad2f33615e56174a1abf6da168cebfa8868f4ba273f16b7, 256'h20aa73ffe48afa6435cd258b173d0c2377d69022e7d098d75caf24c8c5e06b1c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{68, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hfdc70602766f8eed11a6c99a71c973d5659355507b843da6e327a28c11893db9, 256'h3df5349688a085b137b1eacf456a9e9e0f6d15ec0078ca60a7f83f2b10d21350},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{69, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hb516a314f2fce530d6537f6a6c49966c23456f63c643cf8e0dc738f7b876e675, 256'hd39ffd033c92b6d717dd536fbc5efdf1967c4bd80954479ba66b0120cd16fff2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{70, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3b2cbf046eac45842ecb7984d475831582717bebb6492fd0a485c101e29ff0a8, 256'h4c9b7b47a98b0f82de512bc9313aaf51701099cac5f76e68c8595fc1c1d99258},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{71, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h30c87d35e636f540841f14af54e2f9edd79d0312cfa1ab656c3fb15bfde48dcf, 256'h47c15a5a82d24b75c85a692bd6ecafeb71409ede23efd08e0db9abf6340677ed},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{72, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h38686ff0fda2cef6bc43b58cfe6647b9e2e8176d168dec3c68ff262113760f52, 256'h067ec3b651f422669601662167fa8717e976e2db5e6a4cf7c2ddabb3fde9d67d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{73, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h44a3e23bf314f2b344fc25c7f2de8b6af3e17d27f5ee844b225985ab6e2775cf, 256'h2d48e223205e98041ddc87be532abed584f0411f5729500493c9cc3f4dd15e86},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{74, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ded5b7ec8e90e7bf11f967a3d95110c41b99db3b5aa8d330eb9d638781688e9, 256'h7d5792c53628155e1bfc46fb1a67e3088de049c328ae1f44ec69238a009808f9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{75, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hbdae7bcb580bf335efd3bc3d31870f923eaccafcd40ec2f605976f15137d8b8f, 256'hf6dfa12f19e525270b0106eecfe257499f373a4fb318994f24838122ce7ec3c7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{76, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h50f9c4f0cd6940e162720957ffff513799209b78596956d21ece251c2401f1c6, 256'hd7033a0a787d338e889defaaabb106b95a4355e411a59c32aa5167dfab244726},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{77, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hf612820687604fa01906066a378d67540982e29575d019aabe90924ead5c860d, 256'h3f9367702dd7dd4f75ea98afd20e328a1a99f4857b316525328230ce294b0fef},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{78, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h9505e407657d6e8bc93db5da7aa6f5081f61980c1949f56b0f2f507da5782a7a, 256'hc60d31904e3669738ffbeccab6c3656c08e0ed5cb92b3cfa5e7f71784f9c5021},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{79, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hbbd16fbbb656b6d0d83e6a7787cd691b08735aed371732723e1c68a40404517d, 256'h9d8e35dba96028b7787d91315be675877d2d097be5e8ee34560e3e7fd25c0f00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{80, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2ec9760122db98fd06ea76848d35a6da442d2ceef7559a30cf57c61e92df327e, 256'h7ab271da90859479701fccf86e462ee3393fb6814c27b760c4963625c0a19878},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{81, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h54e76b7683b6650baa6a7fc49b1c51eed9ba9dd463221f7a4f1005a89fe00c59, 256'h2ea076886c773eb937ec1cc8374b7915cfd11b1c1ae1166152f2f7806a31c8fd},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{82, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5291deaf24659ffbbce6e3c26f6021097a74abdbb69be4fb10419c0c496c9466, 256'h65d6fcf336d27cc7cdb982bb4e4ecef5827f84742f29f10abf83469270a03dc3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{83, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h207a3241812d75d947419dc58efb05e8003b33fc17eb50f9d15166a88479f107, 256'hcdee749f2e492b213ce80b32d0574f62f1c5d70793cf55e382d5caadf7592767},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{84, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6554e49f82a855204328ac94913bf01bbe84437a355a0a37c0dee3cf81aa7728, 256'haea00de2507ddaf5c94e1e126980d3df16250a2eaebc8be486effe7f22b4f929},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{85, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'ha54c5062648339d2bff06f71c88216c26c6e19b4d80a8c602990ac82707efdfc, 256'he99bbe7fcfafae3e69fd016777517aa01056317f467ad09aff09be73c9731b0d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{86, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h975bd7157a8d363b309f1f444012b1a1d23096593133e71b4ca8b059cff37eaf, 256'h7faa7a28b1c822baa241793f2abc930bd4c69840fe090f2aacc46786bf919622},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{87, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5694a6f84b8f875c276afd2ebcfe4d61de9ec90305afb1357b95b3e0da43885e, 256'h0dffad9ffd0b757d8051dec02ebdf70d8ee2dc5c7870c0823b6ccc7c679cbaa4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{88, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'ha0c30e8026fdb2b4b4968a27d16a6d08f7098f1a98d21620d7454ba9790f1ba6, 256'h5e470453a8a399f15baf463f9deceb53acc5ca64459149688bd2760c65424339},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{89, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h614ea84acf736527dd73602cd4bb4eea1dfebebd5ad8aca52aa0228cf7b99a88, 256'h737cc85f5f2d2f60d1b8183f3ed490e4de14368e96a9482c2a4dd193195c902f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{90, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hbead6734ebe44b810d3fb2ea00b1732945377338febfd439a8d74dfbd0f942fa, 256'h6bb18eae36616a7d3cad35919fd21a8af4bbe7a10f73b3e036a46b103ef56e2a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{91, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h499625479e161dacd4db9d9ce64854c98d922cbf212703e9654fae182df9bad2, 256'h42c177cf37b8193a0131108d97819edd9439936028864ac195b64fca76d9d693},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{92, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h08f16b8093a8fb4d66a2c8065b541b3d31e3bfe694f6b89c50fb1aaa6ff6c9b2, 256'h9d6455e2d5d1779748573b611cb95d4a21f967410399b39b535ba3e5af81ca2e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{93, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hbe26231b6191658a19dd72ddb99ed8f8c579b6938d19bce8eed8dc2b338cb5f8, 256'he1d9a32ee56cffed37f0f22b2dcb57d5c943c14f79694a03b9c5e96952575c89},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{94, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h15e76880898316b16204ac920a02d58045f36a229d4aa4f812638c455abe0443, 256'he74d357d3fcb5c8c5337bd6aba4178b455ca10e226e13f9638196506a1939123},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{95, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h352ecb53f8df2c503a45f9846fc28d1d31e6307d3ddbffc1132315cc07f16dad, 256'h1348dfa9c482c558e1d05c5242ca1c39436726ecd28258b1899792887dd0a3c6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{96, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4a40801a7e606ba78a0da9882ab23c7677b8642349ed3d652c5bfa5f2a9558fb, 256'h3a49b64848d682ef7f605f2832f7384bdc24ed2925825bf8ea77dc5981725782},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{97, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'heacc5e1a8304a74d2be412b078924b3bb3511bac855c05c9e5e9e44df3d61e96, 256'h7451cd8e18d6ed1885dd827714847f96ec4bb0ed4c36ce9808db8f714204f6d1},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{98, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2f7a5e9e5771d424f30f67fdab61e8ce4f8cd1214882adb65f7de94c31577052, 256'hac4e69808345809b44acb0b2bd889175fb75dd050c5a449ab9528f8f78daa10c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{99, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffcda40f792ce4d93e7e0f0e95e1a2147dddd7f6487621c30a03d710b3300219, 256'h79938b55f8a17f7ed7ba9ade8f2065a1fa77618f0b67add8d58c422c2453a49a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{100, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h81f2359c4faba6b53d3e8c8c3fcc16a948350f7ab3a588b28c17603a431e39a8, 256'hcd6f6a5cc3b55ead0ff695d06c6860b509e46d99fccefb9f7f9e101857f74300},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{101, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdfc8bf520445cbb8ee1596fb073ea283ea130251a6fdffa5c3f5f2aaf75ca808, 256'h048e33efce147c9dd92823640e338e68bfd7d0dc7a4905b3a7ac711e577e90e7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{102, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'had019f74c6941d20efda70b46c53db166503a0e393e932f688227688ba6a5762, 256'h93320eb7ca0710255346bdbb3102cdcf7964ef2e0988e712bc05efe16c199345},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{103, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hac8096842e8add68c34e78ce11dd71e4b54316bd3ebf7fffdeb7bd5a3ebc1883, 256'hf5ca2f4f23d674502d4caf85d187215d36e3ce9f0ce219709f21a3aac003b7a8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{104, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h677b2d3a59b18a5ff939b70ea002250889ddcd7b7b9d776854b4943693fb92f7, 256'h6b4ba856ade7677bf30307b21f3ccda35d2f63aee81efd0bab6972cc0795db55},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{105, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h479e1ded14bcaed0379ba8e1b73d3115d84d31d4b7c30e1f05e1fc0d5957cfb0, 256'h918f79e35b3d89487cf634a4f05b2e0c30857ca879f97c771e877027355b2443},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{106, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h43dfccd0edb9e280d9a58f01164d55c3d711e14b12ac5cf3b64840ead512a0a3, 256'h1dbe33fa8ba84533cd5c4934365b3442ca1174899b78ef9a3199f49584389772},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{107, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5b09ab637bd4caf0f4c7c7e4bca592fea20e9087c259d26a38bb4085f0bbff11, 256'h45b7eb467b6748af618e9d80d6fdcd6aa24964e5a13f885bca8101de08eb0d75},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{108, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5e9b1c5a028070df5728c5c8af9b74e0667afa570a6cfa0114a5039ed15ee06f, 256'hb1360907e2d9785ead362bb8d7bd661b6c29eeffd3c5037744edaeb9ad990c20},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{109, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0671a0a85c2b72d54a2fb0990e34538b4890050f5a5712f6d1a7a5fb8578f32e, 256'hdb1846bab6b7361479ab9c3285ca41291808f27fd5bd4fdac720e5854713694c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{110, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7673f8526748446477dbbb0590a45492c5d7d69859d301abbaedb35b2095103a, 256'h3dc70ddf9c6b524d886bed9e6af02e0e4dec0d417a414fed3807ef4422913d7c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{111, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7f085441070ecd2bb21285089ebb1aa6450d1a06c36d3ff39dfd657a796d12b5, 256'h249712012029870a2459d18d47da9aa492a5e6cb4b2d8dafa9e4c5c54a2b9a8b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{112, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h914c67fb61dd1e27c867398ea7322d5ab76df04bc5aa6683a8e0f30a5d287348, 256'hfa07474031481dda4953e3ac1959ee8cea7e66ec412b38d6c96d28f6d37304ea},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{113, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0ad99500288d466940031d72a9f5445a4d43784640855bf0a69874d2de5fe103, 264'h00c5011e6ef2c42dcd50d5d3d29f99ae6eba2c80c9244f4c5422f0979ff0c3ba5e, 256'h000000000000000000000000000000004319055358e8617b0c46353d039cdaab, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{114, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0ad99500288d466940031d72a9f5445a4d43784640855bf0a69874d2de5fe103, 264'h00c5011e6ef2c42dcd50d5d3d29f99ae6eba2c80c9244f4c5422f0979ff0c3ba5e, 256'hffffffff00000001000000000000000000000000fffffffffffffffffffffffc, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{115, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00ab05fd9d0de26b9ce6f4819652d9fc69193d0aa398f0fba8013e09c582204554, 256'h19235271228c786759095d12b75af0692dd4103f19f6a8c32f49435a1e9b8d45, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254f, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{116, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0080984f39a1ff38a86a68aa4201b6be5dfbfecf876219710b07badf6fdd4c6c56, 256'h11feb97390d9826e7a06dfb41871c940d74415ed3cac2089f1445019bb55ed95, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h909135bdb6799286170f5ead2de4f6511453fe50914f3df2de54a36383df8dd4},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{117, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4201b4272944201c3294f5baa9a3232b6dd687495fcc19a70a95bc602b4f7c05, 264'h0095c37eba9ee8171c1bb5ac6feaf753bc36f463e3aef16629572c0c0a8fb0800e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h27b4577ca009376f71303fd5dd227dcef5deb773ad5f5a84360644669ca249a5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{118, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a71af64de5126a4a4e02b7922d66ce9415ce88a4c9d25514d91082c8725ac957, 256'h5d47723c8fbe580bb369fec9c2665d8e30a435b9932645482e7c9f11e872296b, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{119, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a71af64de5126a4a4e02b7922d66ce9415ce88a4c9d25514d91082c8725ac957, 256'h5d47723c8fbe580bb369fec9c2665d8e30a435b9932645482e7c9f11e872296b, 8'h05, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{120, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6627cec4f0731ea23fc2931f90ebe5b7572f597d20df08fc2b31ee8ef16b1572, 256'h6170ed77d8d0a14fc5c9c3c4c9be7f0d3ee18f709bb275eaf2073e258fe694a5, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000003},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{121, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6627cec4f0731ea23fc2931f90ebe5b7572f597d20df08fc2b31ee8ef16b1572, 256'h6170ed77d8d0a14fc5c9c3c4c9be7f0d3ee18f709bb275eaf2073e258fe694a5, 8'h05, 8'h03},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{122, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5a7c8825e85691cce1f5e7544c54e73f14afc010cb731343262ca7ec5a77f5bf, 264'h00ef6edf62a4497c1bd7b147fb6c3d22af3c39bfce95f30e13a16d3d7b2812f813, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000005},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{123, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5a7c8825e85691cce1f5e7544c54e73f14afc010cb731343262ca7ec5a77f5bf, 264'h00ef6edf62a4497c1bd7b147fb6c3d22af3c39bfce95f30e13a16d3d7b2812f813, 8'h05, 8'h05},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{124, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00cbe0c29132cd738364fedd603152990c048e5e2fff996d883fa6caca7978c737, 256'h70af6a8ce44cb41224b2603606f4c04d188e80bff7cc31ad5189d4ab0d70e8c1, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000006},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{125, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00cbe0c29132cd738364fedd603152990c048e5e2fff996d883fa6caca7978c737, 256'h70af6a8ce44cb41224b2603606f4c04d188e80bff7cc31ad5189d4ab0d70e8c1, 8'h05, 8'h06},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00cbe0c29132cd738364fedd603152990c048e5e2fff996d883fa6caca7978c737, 256'h70af6a8ce44cb41224b2603606f4c04d188e80bff7cc31ad5189d4ab0d70e8c1, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632556, 256'h0000000000000000000000000000000000000000000000000000000000000006},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4be4178097002f0deab68f0d9a130e0ed33a6795d02a20796db83444b037e139, 256'h20f13051e0eecdcfce4dacea0f50d1f247caa669f193c1b4075b51ae296d2d56, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc75fbd8},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{128, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d0f73792203716afd4be4329faa48d269f15313ebbba379d7783c97bf3e890d9, 264'h00971f4a3206605bec21782bf5e275c714417e8f566549e6bc68690d2363c89cc1, 256'h0000000000000000000000000000000000000000000000000000000000000100, 256'h8f1e3c7862c58b16bb76eddbb76eddbb516af4f63f2d74d76e0d28c9bb75ea88},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{129, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4838b2be35a6276a80ef9e228140f9d9b96ce83b7a254f71ccdebbb8054ce05f, 264'h00fa9cbc123c919b19e00238198d04069043bd660a828814051fcb8aac738a6c6b, 256'h000000000000000000000000000000000000000000000000002d9b4d347952d6, 256'hef3043e7329581dbb3974497710ab11505ee1c87ff907beebadd195a0ffe6d7a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{130, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h7393983ca30a520bbc4783dc9960746aab444ef520c0a8e771119aa4e74b0f64, 264'h00e9d7be1ab01a0bf626e709863e6a486dbaf32793afccf774e2c6cd27b1857526, 256'h000000000000000000000000000000000000001033e67e37b32b445580bf4eff, 256'h8b748b74000000008b748b748b748b7466e769ad4a16d3dcd87129b8e91d1b4d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{131, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5ac331a1103fe966697379f356a937f350588a05477e308851b8a502d5dfcdc5, 264'h00fe9993df4b57939b2b8da095bf6d794265204cfe03be995a02e65d408c871c0b, 256'h0000000000000000000000000000000000000000000000000000000000000100, 256'hef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{132, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1d209be8de2de877095a399d3904c74cc458d926e27bb8e58e5eae5767c41509, 264'h00dd59e04c214f7b18dce351fc2a549893a6860e80163f38cc60a4f2c9d040d8c9, 256'h00000000000000000000000000000000000000062522bbd3ecbe7c39e93e7c25, 256'hef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{133, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h083539fbee44625e3acaafa2fcb41349392cef0633a1b8fabecee0c133b10e99, 264'h00915c1ebe7bf00df8535196770a58047ae2a402f26326bb7d41d4d7616337911e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc6324d5, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{134, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008aeb368a7027a4d64abdea37390c0c1d6a26f399e2d9734de1eb3d0e19373874, 256'h05bd13834715e1dbae9b875cf07bd55e1b6691c7f7536aef3b19bf7a4adf576d, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008aeb368a7027a4d64abdea37390c0c1d6a26f399e2d9734de1eb3d0e19373874, 256'h05bd13834715e1dbae9b875cf07bd55e1b6691c7f7536aef3b19bf7a4adf576d, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{136, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b533d4695dd5b8c5e07757e55e6e516f7e2c88fa0239e23f60e8ec07dd70f287, 256'h1b134ee58cc583278456863f33c3a85d881f7d4a39850143e29d4eaf009afe47, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{137, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f50d371b91bfb1d7d14e1323523bc3aa8cbf2c57f9e284de628c8b4536787b86, 264'h00f94ad887ac94d527247cd2e7d0c8b1291c553c9730405380b14cbb209f5fa2dd, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{138, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h68ec6e298eafe16539156ce57a14b04a7047c221bafc3a582eaeb0d857c4d946, 264'h0097bed1af17850117fdb39b2324f220a5698ed16c426a27335bb385ac8ca6fb30, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{139, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h69da0364734d2e530fece94019265fefb781a0f1b08f6c8897bdf6557927c8b8, 256'h66d2d3c7dcd518b23d726960f069ad71a933d86ef8abbcce8b20f71e2a847002, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{140, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d8adc00023a8edc02576e2b63e3e30621a471e2b2320620187bf067a1ac1ff32, 256'h33e2b50ec09807accb36131fff95ed12a09a86b4ea9690aa32861576ba2362e1, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h44a5ad0ad0636d9f12bc9e0a6bdd5e1cbcb012ea7bf091fcec15b0c43202d52e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{141, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3623ac973ced0a56fa6d882f03a7d5c7edca02cfc7b2401fab3690dbe75ab785, 264'h008db06908e64b28613da7257e737f39793da8e713ba0643b92e9bb3252be7f8fe, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{142, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00cf04ea77e9622523d894b93ff52dc3027b31959503b6fa3890e5e04263f922f1, 264'h00e8528fb7c006b3983c8b8400e57b4ed71740c2f3975438821199bedeaecab2e9, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'haaaaaaaa00000000aaaaaaaaaaaaaaaa7def51c91a0fbf034d26872ca84218e1},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{143, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00db7a2c8a1ab573e5929dc24077b508d7e683d49227996bda3e9f78dbeff77350, 256'h4f417f3bc9a88075c2e0aadd5a13311730cf7cc76a82f11a36eaf08a6c99a206, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'he91e1ba60fdedb76a46bcb51dc0b8b4b7e019f0a28721885fa5d3a8196623397},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{144, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00dead11c7a5b396862f21974dc4752fadeff994efe9bbd05ab413765ea80b6e1f, 256'h1de3f0640e8ac6edcf89cff53c40e265bb94078a343736df07aa0318fc7fe1ff, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hfdea5843ffeb73af94313ba4831b53fe24f799e525b1e8e8c87b59b95b430ad9},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{145, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d0bc472e0d7c81ebaed3a6ef96c18613bb1fea6f994326fbe80e00dfde67c7e9, 264'h00986c723ea4843d48389b946f64ad56c83ad70ff17ba85335667d1bb9fa619efd, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h03ffcabf2f1b4d2a65190db1680d62bb994e41c5251cd73b3c3dfc5e5bafc035},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{146, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a0a44ca947d66a2acb736008b9c08d1ab2ad03776e02640f78495d458dd51c32, 256'h6337fe5cf8c4604b1f1c409dc2d872d4294a4762420df43a30a2392e40426add, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h4dfbc401f971cd304b33dfdb17d0fed0fe4c1a88ae648e0d2847f74977534989},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{147, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00c9c2115290d008b45fb65fad0f602389298c25420b775019d42b62c3ce8a96b7, 256'h3877d25a8080dc02d987ca730f0405c2c9dbefac46f9e601cc3f06e9713973fd, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbc4024761cd2ffd43dfdb17d0fed112b988977055cd3a8e54971eba9cda5ca71},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{148, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5eca1ef4c287dddc66b8bccf1b88e8a24c0018962f3c5e7efa83bc1a5ff6033e, 256'h5e79c4cb2c245b8c45abdce8a8e4da758d92a607c32cd407ecaef22f1c934a71, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h788048ed39a5ffa77bfb62fa1fda2257742bf35d128fb3459f2a0c909ee86f91},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{149, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5caaa030e7fdf0e4936bc7ab5a96353e0a01e4130c3f8bf22d473e317029a47a, 264'h00deb6adc462f7058f2a20d371e9702254e9b201642005b3ceda926b42b178bef9, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h476d9131fd381bd917d0fed112bc9e0a5924b5ed5b11167edd8b23582b3cb15e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{150, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00c2fd20bac06e555bb8ac0ce69eb1ea20f83a1fc3501c8a66469b1a31f619b098, 256'h6237050779f52b615bd7b8d76a25fc95ca2ed32525c75f27ffc87ac397e6cbaf, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h8374253e3e21bd154448d0a8f640fe46fafa8b19ce78d538f6cc0a19662d3601},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{151, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3fd6a1ca7f77fb3b0bbe726c372010068426e11ea6ae78ce17bedae4bba86ced, 256'h03ce5516406bf8cfaab8745eac1cd69018ad6f50b5461872ddfc56e0db3c8ff4, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h357cfd3be4d01d413c5b9ede36cba5452c11ee7fe14879e749ae6a2d897a52d6},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{152, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h009cb8e51e27a5ae3b624a60d6dc32734e4989db20e9bca3ede1edf7b086911114, 264'h00b4c104ab3c677e4b36d6556e8ad5f523410a19f2e277aa895fc57322b4427544, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h29798c5c0ee287d4a5e8e6b799fd86b8df5225298e6ffc807cd2f2bc27a0a6d8},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{153, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a3e52c156dcaf10502620b7955bc2b40bc78ef3d569e1223c262512d8f49602a, 256'h4a2039f31c1097024ad3cc86e57321de032355463486164cf192944977df147f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h0b70f22c781092452dca1a5711fa3a5a1f72add1bf52c2ff7cae4820b30078dd},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{154, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f19b78928720d5bee8e670fb90010fb15c37bf91b58a5157c3f3c059b2655e88, 264'h00cf701ec962fb4a11dcf273f5dc357e58468560c7cfeb942d074abd4329260509, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h16e1e458f021248a5b9434ae23f474b43ee55ba37ea585fef95c90416600f1ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{155, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0083a744459ecdfb01a5cf52b27a05bb7337482d242f235d7b4cb89345545c90a8, 264'h00c05d49337b9649813287de9ffe90355fd905df5f3c32945828121f37cc50de6e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h2252d6856831b6cf895e4f0535eeaf0e5e5809753df848fe760ad86219016a97},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{156, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00dd13c6b34c56982ddae124f039dfd23f4b19bbe88cee8e528ae51e5d6f3a21d7, 264'h00bfad4c2e6f263fe5eb59ca974d039fc0e4c3345692fb5320bdae4bd3b42a45ff, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h81ffe55f178da695b28c86d8b406b15dab1a9e39661a3ae017fbe390ac0972c3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{157, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h67e6f659cdde869a2f65f094e94e5b4dfad636bbf95192feeed01b0f3deb7460, 264'h00a37e0a51f258b7aeb51dfe592f5cfd5685bbe58712c8d9233c62886437c38ba0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffffaaaaaaaaffffffffffffffffe9a2538f37b28a2c513dee40fecbb71a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{158, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2eb6412505aec05c6545f029932087e490d05511e8ec1f599617bb367f9ecaaf, 264'h00805f51efcc4803403f9b1ae0124890f06a43fedcddb31830f6669af292895cb0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hb62f26b5f2a2b26f6de86d42ad8a13da3ab3cccd0459b201de009e526adf21f2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{159, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0084db645868eab35e3a9fd80e056e2e855435e3a6b68d75a50a854625fe0d7f35, 256'h6d2589ac655edc9a11ef3e075eddda9abf92e72171570ef7bf43a2ee39338cfe, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbb1d9ac949dd748cd02bbbe749bd351cd57b38bb61403d700686aa7b4c90851e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{160, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0091b9e47c56278662d75c0983b22ca8ea6aa5059b7a2ff7637eb2975e386ad663, 256'h49aa8ff283d0f77c18d6d11dc062165fd13c3c0310679c1408302a16854ecfbd, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h66755a00638cdaec1c732513ca0234ece52545dac11f816e818f725b4f60aaf2},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{161, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f3ec2f13caf04d0192b47fb4c5311fb6d4dc6b0a9e802e5327f7ec5ee8e4834d, 264'h00f97e3e468b7d0db867d6ecfe81e2b0f9531df87efdb47c1338ac321fefe5a432, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h55a00c9fcdaebb6032513ca0234ecfffe98ebe492fdf02e48ca48e982beb3669},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{162, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d92b200aefcab6ac7dafd9acaf2fa10b3180235b8f46b4503e4693c670fccc88, 256'h5ef2f3aebf5b317475336256768f7c19efb7352d27e4cccadc85b6b8ab922c72, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hab40193f9b5d76c064a27940469d9fffd31d7c925fbe05c919491d3057d66cd2},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{163, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0a88361eb92ecca2625b38e5f98bbabb96bf179b3d76fc48140a3bcd881523cd, 264'h00e6bdf56033f84a5054035597375d90866aa2c96b86a41ccf6edebf47298ad489, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hca0234ebb5fdcb13ca0234ecffffffffcb0dadbbc7f549f8a26b4408d0dc8600},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{164, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d0fb17ccd8fafe827e0c1afc5d8d80366e2b20e7f14a563a2ba50469d84375e8, 256'h68612569d39e2bb9f554355564646de99ac602cc6349cf8c1e236a7de7637d93, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbfffffff3ea3677e082b9310572620ae19933a9e65b285598711c77298815ad3},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{165, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00836f33bbc1dc0d3d3abbcef0d91f11e2ac4181076c9af0a22b1e4309d3edb276, 264'h009ab443ff6f901e30c773867582997c2bec2b0cb8120d760236f3a95bbe881f75, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h266666663bbbbbbbe6666666666666665b37902e023fab7c8f055d86e5cc41f4},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{166, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0092f99fbe973ed4a299719baee4b432741237034dec8d72ba5103cb33e55feeb8, 256'h033dd0e91134c734174889f3ebcf1b7a1ac05767289280ee7a794cebd6e69697, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbfffffff36db6db7a492492492492492146c573f4c6dfc8d08a443e258970b09},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{167, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d35ba58da30197d378e618ec0fa7e2e2d12cffd73ebbb2049d130bba434af09e, 264'h00ff83986e6875e41ea432b7585a49b3a6c77cbb3c47919f8e82874c794635c1d2, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbfffffff2aaaaaab7fffffffffffffffc815d0e60b3e596ecb1ad3a27cfd49c4},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{168, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008651ce490f1b46d73f3ff475149be29136697334a519d7ddab0725c8d0793224, 264'h00e11c65bd8ca92dc8bc9ae82911f0b52751ce21dd9003ae60900bd825f590cc28, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffff55555555ffffffffffffffffd344a71e6f651458a27bdc81fd976e37},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{169, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6d8e1b12c831a0da8795650ff95f101ed921d9e2f72b15b1cdaca9826b9cfc6d, 264'h00ef6d63e2bc5c089570394a4bc9f892d5e6c7a6a637b20469a58c106ad486bf37, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h3fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192aa},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{170, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0ae580bae933b4ef2997cbdbb0922328ca9a410f627a0f7dff24cb4d920e1542, 264'h008911e7f8cc365a8a88eb81421a361ccc2b99e309d8dcd9a98ba83c3949d893e3, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5d8ecd64a4eeba466815ddf3a4de9a8e6abd9c5db0a01eb80343553da648428f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{171, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5b812fd521aafa69835a849cce6fbdeb6983b442d2444fe70e134c027fc46963, 264'h00838a40f2a36092e9004e92d8d940cf5638550ce672ce8b8d4e15eba5499249e9, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 256'hbb726660235793aa9957a61e76e00c2c435109cf9a15dd624d53f4301047856b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5b812fd521aafa69835a849cce6fbdeb6983b442d2444fe70e134c027fc46963, 256'h7c75bf0c5c9f6d17ffb16d2726bf30a9c7aaf31a8d317472b1ea145ab66db616, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 256'hbb726660235793aa9957a61e76e00c2c435109cf9a15dd624d53f4301047856b},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6adda82b90261b0f319faa0d878665a6b6da497f09c903176222c34acfef72a6, 256'h47e6f50dcc40ad5d9b59f7602bb222fad71a41bf5e1f9df4959a364c62e488d9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00dd86d3b5f4a13e8511083b78002081c53ff467f11ebd98a51a633db76665d250, 256'h45d5c8200c89f2fa10d849349226d21d8dfaed6ff8d5cb3e1b7e17474ebc18f7, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{176, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4fea55b32cb32aca0c12c4cd0abfb4e64b0f5a516e578c016591a93f5a0fbcc5, 264'h00d7d3fd10b2be668c547b212f6bb14c88f0fecd38a8a4b2c785ed3be62ce4b280, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{177, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00c6a771527024227792170a6f8eee735bf32b7f98af669ead299802e32d7c3107, 264'h00bc3b4b5e65ab887bbd343572b3e5619261fe3a073e2ffd78412f726867db589e, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'hb6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{178, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00851c2bbad08e54ec7a9af99f49f03644d6ec6d59b207fec98de85a7d15b956ef, 264'h00cee9960283045075684b410be8d0f7494b91aa2379f60727319f10ddeb0fe9d6, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'hcccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{179, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f6417c8a670584e388676949e53da7fc55911ff68318d1bf3061205acb19c48f, 264'h008f2b743df34ad0f72674acb7505929784779cd9ac916c3669ead43026ab6d43f, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{180, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h501421277be45a5eefec6c639930d636032565af420cf3373f557faa7f8a0643, 264'h008673d6cb6076e1cfcdc7dfe7384c8e5cac08d74501f2ae6e89cad195d0aa1371, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{181, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0d935bf9ffc115a527735f729ca8a4ca23ee01a4894adf0e3415ac84e808bb34, 256'h3195a3762fea29ed38912bd9ea6c4fde70c3050893a4375850ce61d82eba33c5, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{182, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5e59f50708646be8a589355014308e60b668fb670196206c41e748e64e4dca21, 256'h5de37fee5c97bcaf7144d5b459982f52eeeafbdf03aacbafef38e213624a01de, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{183, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h169fb797325843faff2f7a5b5445da9e2fd6226f7ef90ef0bfe924104b02db8e, 256'h7bbb8de662c7b9b1cf9b22f7a2e582bd46d581d68878efb2b861b131d8a1d667, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'hb6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{184, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h271cd89c000143096b62d4e9e4ca885aef2f7023d18affdaf8b7b54898148754, 256'h0a1c6e954e32108435b55fa385b0f76481a609b9149ccb4b02b2ca47fe8e4da5, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'hcccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{185, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3d0bc7ed8f09d2cb7ddb46ebc1ed799ab1563a9ab84bf524587a220afe499c12, 264'h00e22dc3b3c103824a4f378d96adb0a408abf19ce7d68aa6244f78cb216fa3f8df, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{186, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a6c885ade1a4c566f9bb010d066974abb281797fa701288c721bcbd23663a9b7, 256'h2e424b690957168d193a6096fc77a2b004a9c7d467e007e1f2058458f98af316, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{187, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008d3c2c2c3b765ba8289e6ac3812572a25bf75df62d87ab7330c3bdbad9ebfa5c, 256'h4c6845442d66935b238578d43aec54f7caa1621d1af241d4632e0b780c423f5d, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{188, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{189, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'h44a5ad0ad0636d9f12bc9e0a6bdd5e1cbcb012ea7bf091fcec15b0c43202d52e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{190, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'h44a5ad0ad0636d9f12bc9e0a6bdd5e1cbcb012ea7bf091fcec15b0c43202d52e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{192, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'hb292a619339f6e567a305c951c0dcbcc42d16e47f219f9e98e76e09d8770b34a, 256'h0177e60492c5a8242f76f07bfe3661bde59ec2a17ce5bd2dab2abebdf89a62e2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{193, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h530bd6b0c9af2d69ba897f6b5fb59695cfbf33afe66dbadcf5b8d2a2a6538e23, 256'hd85e489cb7a161fd55ededcedbf4cc0c0987e3e3f0f242cae934c72caa3f43e9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{194, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'ha8ea150cb80125d7381c4c1f1da8e9de2711f9917060406a73d7904519e51388, 256'hf3ab9fa68bd47973a73b2d40480c2ba50c22c9d76ec217257288293285449b86},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{195, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h986e65933ef2ed4ee5aada139f52b70539aaf63f00a91f29c69178490d57fb71, 256'h3dafedfb8da6189d372308cbf1489bbbdabf0c0217d1c0ff0f701aaa7a694b9c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{196, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'hd434e262a49eab7781e353a3565e482550dd0fd5defa013c7f29745eff3569f1, 256'h9b0c0a93f267fb6052fd8077be769c2b98953195d7bc10de844218305c6ba17a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{197, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h0fe774355c04d060f76d79fd7a772e421463489221bf0a33add0be9b1979110b, 256'h500dcba1c69a8fbd43fa4f57f743ce124ca8b91a1f325f3fac6181175df55737},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{198, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'hbb40bf217bed3fb3950c7d39f03d36dc8e3b2cd79693f125bfd06595ee1135e3, 256'h541bf3532351ebb032710bdb6a1bf1bfc89a1e291ac692b3fa4780745bb55677},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{199, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h664eb7ee6db84a34df3c86ea31389a5405badd5ca99231ff556d3e75a233e73a, 256'h59f3c752e52eca46137642490a51560ce0badc678754b8f72e51a2901426a1bd},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{200, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h4cd0429bbabd2827009d6fcd843d4ce39c3e42e2d1631fd001985a79d1fd8b43, 256'h9638bf12dd682f60be7ef1d0e0d98f08b7bca77a1a2b869ae466189d2acdabe3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{201, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'he56c6ea2d1b017091c44d8b6cb62b9f460e3ce9aed5e5fd41e8added97c56c04, 256'ha308ec31f281e955be20b457e463440b4fcf2b80258078207fc1378180f89b55},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{202, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h1158a08d291500b4cabed3346d891eee57c176356a2624fb011f8fbbf3466830, 256'h228a8c486a736006e082325b85290c5bc91f378b75d487dda46798c18f285519},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{203, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'hb1db9289649f59410ea36b0c0fc8d6aa2687b29176939dd23e0dde56d309fa9d, 256'h3e1535e4280559015b0dbd987366dcf43a6d1af5c23c7d584e1c3f48a1251336},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{204, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'hb7b16e762286cb96446aa8d4e6e7578b0a341a79f2dd1a220ac6f0ca4e24ed86, 256'hddc60a700a139b04661c547d07bbb0721780146df799ccf55e55234ecb8f12bc},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{205, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'hd82a7c2717261187c8e00d8df963ff35d796edad36bc6e6bd1c91c670d9105b4, 256'h3dcabddaf8fcaa61f4603e7cbac0f3c0351ecd5988efb23f680d07debd139929},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{206, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'h5eb9c8845de68eb13d5befe719f462d77787802baff30ce96a5cba063254af78, 256'h2c026ae9be2e2a5e7ca0ff9bbd92fb6e44972186228ee9a62b87ddbe2ef66fb5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{207, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'h96843dd03c22abd2f3b782b170239f90f277921becc117d0404a8e4e36230c28, 256'hf2be378f526f74a543f67165976de9ed9a31214eb4d7e6db19e1ede123dd991d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{208, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h766456dce1857c906f9996af729339464d27e9d98edc2d0e3b760297067421f6, 256'h402385ecadae0d8081dccaf5d19037ec4e55376eced699e93646bfbbf19d0b41},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{209, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'hc605c4b2edeab20419e6518a11b2dbc2b97ed8b07cced0b19c34f777de7b9fd9, 256'hedf0f612c5f46e03c719647bc8af1b29b2cde2eda700fb1cff5e159d47326dba},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{210, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'hd48b68e6cabfe03cf6141c9ac54141f210e64485d9929ad7b732bfe3b7eb8a84, 256'hfeedae50c61bd00e19dc26f9b7e2265e4508c389109ad2f208f0772315b6c941},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{211, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'hb7c81457d4aeb6aa65957098569f0479710ad7f6595d5874c35a93d12a5dd4c7, 256'hb7961a0b652878c2d568069a432ca18a1a9199f2ca574dad4b9e3a05c0a1cdb3},  // lens: hash=256b(32B), x=232b(29B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{212, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h6b01332ddb6edfa9a30a1321d5858e1ee3cf97e263e669f8de5e9652e76ff3f7, 256'h5939545fced457309a6a04ace2bd0f70139c8f7d86b02cb1cc58f9e69e96cd5a},  // lens: hash=256b(32B), x=232b(29B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{213, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'hefdb884720eaeadc349f9fc356b6c0344101cd2fd8436b7d0e6a4fb93f106361, 256'hf24bee6ad5dc05f7613975473aadf3aacba9e77de7d69b6ce48cb60d8113385d},  // lens: hash=256b(32B), x=232b(29B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{214, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h31230428405560dcb88fb5a646836aea9b23a23dd973dcbe8014c87b8b20eb07, 256'h0f9344d6e812ce166646747694a41b0aaf97374e19f3c5fb8bd7ae3d9bd0beff},  // lens: hash=256b(32B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{215, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'hcaa797da65b320ab0d5c470cda0b36b294359c7db9841d679174db34c4855743, 256'hcf543a62f23e212745391aaf7505f345123d2685ee3b941d3de6d9b36242e5a0},  // lens: hash=256b(32B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{216, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h7e5f0ab5d900d3d3d7867657e5d6d36519bc54084536e7d21c336ed800185945, 256'h9450c07f201faec94b82dfb322e5ac676688294aad35aa72e727ff0b19b646aa},  // lens: hash=256b(32B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{217, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'hd7d70c581ae9e3f66dc6a480bf037ae23f8a1e4a2136fe4b03aa69f0ca25b356, 256'h89c460f8a5a5c2bbba962c8a3ee833a413e85658e62a59e2af41d9127cc47224},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{218, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h341c1b9ff3c83dd5e0dfa0bf68bcdf4bb7aa20c625975e5eeee34bb396266b34, 256'h72b69f061b750fd5121b22b11366fad549c634e77765a017902a67099e0a4469},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{219, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h70bebe684cdcb5ca72a42f0d873879359bd1781a591809947628d313a3814f67, 256'haec03aca8f5587a4d535fa31027bbe9cc0e464b1c3577f4c2dcde6b2094798a9}  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
};
`endif // WYCHERPROOF_SECP256R1_SHA256_P1363_SV
