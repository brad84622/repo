`ifndef WYCHERPROOF_SECP224R1_SHA512_SV
`define WYCHERPROOF_SECP224R1_SHA512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224r1_sha512;

localparam int TEST_VECTORS_SECP224R1_SHA512_NUM = 88;

ecdsa_vector_secp224r1_sha512 test_vectors_secp224r1_sha512 [] = '{
  '{1, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'h394766fb67a65fe0af6c154f7cbd285ea180b4c6150cdafafb0f6f0f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{2, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'hc6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{115, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=0b(0B)
  '{124, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{130, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{139, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'hc6b899049859a01f5093eab08342d7a15e7f4b39eaf3250504f090f1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{143, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'h394766fb67a65fe0af6c154f7cbe11bbc0c7c488012fb1b59eb344d2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{144, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{230, 1'b1, 512'hf582f7e1597d4966b5873f6fb0211f38c289b14924aa3830aa767732dbda99f309d9c9561dcb6255ac12355838d8587b8bb0d09d5f693189904337c73ee68378, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 224'h221a25eb9cc8dd66fdf156b2f6ab601ab6d9c509247f8de5d2671a96},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{231, 1'b1, 512'h0000000001b99889c891f2468c618149cb6865b933cca31eddb353de09746b540616ba69c5f5ff992c6d6177427daf1cb46a4c5c08625263a615fbf3eeaae178, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3b3008ed596b7fa276498def40d96b1eb2ffb731a44050ffb732e4e6, 224'h6dbb08c56db737e9392ff4f3a54d8b806d70af226ecf413b3465de55},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{236, 1'b1, 512'hef200f1a5400000000399e032faaf4b3c32d804555abf20471a3a18dc46f3917eb9072220b5d5f994d27b221346631c47eb579d69cc5e438b7e7b963bca9d84f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7fd45528eb7bfc3710e273c4468f0b50ebf93f94cd0e7a602a4929a6, 224'h46613dd1ffd85df8d71f3498001721fda4982c27a1c291359b05b1b8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{239, 1'b1, 512'hd40c1a66696b7a6500000000ebb22b0b1f80b394770ad61c5c42ff0584ed4c84a3d185d3c07725f0d3080b451dad86945cc9b0801c01e0b6b8739ff8ec36df22, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4314a2bd139d47be3d9fd9ebdd72a06a220219c7596b944178ee6f5f, 224'h0e6f1d2f57c699654e9c705d7b8fa3c1ccb0f939f6368bed246b2e10},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{241, 1'b1, 512'hcf9bb31b573fa12e7e51000000004b37d8761e5d50f214b30bc2b134bc7e0e30653b8debc737a21392357313d13e08eecfdefd8d37bec92b680a84f5430fb57c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h476aaa58677d9e60477cffd026c43248e2cf3cc21e8fdccb75ceefad, 224'h7799fc7af8f9b929203faf899bb5ca1aecf2492555157282dfde790d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{251, 1'b1, 512'hdf8f102f7c54ce2cb6ca609ce724818f7621cdc600000000c69bb15b7c33f6b27c75a153b581d47b99de18ccc8105fc3bb697f180112706c5ebfd6fc6c8a6322, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h785ac8c956d7797ae67498775b3c446c41735eb15f3430b49f6a09f2, 224'h5710879ab83994e809c8d2cbd6f2ac5c205b4b8d6226e98be03e7967},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{256, 1'b1, 512'h295422dc27dfac13c79d2028d3daed64c1dcaad525dbbf14a9000000003667b1baf41fd9137fa0bd8c3851590b206aefb6cde62fb4ecc23ae308e540e83a7f09, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h52a010a23e4f9ebb459bbe9f3057e6c19761fb99d25c9b16b8f007d8, 224'h526dc1f34444de00447ba23c76950f2c159579d548b6335d127ea321},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{259, 1'b1, 512'h057d7524efbce651b92e0a70e4454156e7cd4b696c197c6a064032c100000000768565d4af2019fe3247dba91948292af777f107fdc9c3b47659eaeab26ead77, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1895e65593d71e5635cce022dda19bd155bb9a7f2e307e5ce9127ade, 224'h121b487c320c544dcdd471d46fcde2ce5dc9d17fda70544c4eab50a2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{261, 1'b1, 512'hc7b70cc4a55d55342487a4469ad2243ef6d6b69f11604b8c12baa03dd3e10000000014df0db29a9d4d54b26f4047f3e0c739f7a260768b20589254e1235fc590, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h07a57197667a0c40423d4811ff96384c9330467e8a28eaa4c0d519f4, 224'h011062c8694494baaed24ff610e1e4227efb59a163c33fafd40100f9},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{264, 1'b1, 512'hc0891fc626ef4b106fc00f5c067253f26a2868d09aa2ce029466f353ba525e757100000000a3cee37421995445fae741697659a406394c870d8bdda130080d15, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h596b74077801db2e889d3b2aaa3990fe180abc152d48528385ca955d, 224'h38bffd416f779843fad389750003eb0708112a4834c554f476a3e0d1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{267, 1'b1, 512'hd34ac40ed5ab79a4e5ac1e4081e0e47e4fdedac1555b01ab62a13ac0ae9dbc3c23f799510000000010116f328ad1db0cd68cd1db9e1b34b5a52ebe9b8e372b78, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0a530530b6a9238d2d1a3cf468986c87f3b208f61ea0486d53140c17, 224'h5f027a73f31a5cc2bee81ff0019477c542fd782ecde0e551fcd37e93},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{274, 1'b1, 512'hf1d6ef224f72b83a109944afbfb34ae1f70d6e50eee54a91faf8ba0fc062563113d988f2b826c055ecc61e00000000554878a7e761e75fdf1ed2ad2d138b2974, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h78850a40530aa258e478e7c547d3a5e4944d3524f1676443e4dfb37d, 224'h687058e1ca478f52a30c9a3f8e2eea9d8c40599cd47ef66b9430d17d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{275, 1'b1, 512'hb33f308c5b107050cb2e513fabf8b896e52c85852fbe32308bee8b8661121bdac78f52f924cf3d5690ac92d5000000004f0f619e72ec1464166078ba3f508a66, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h066e7268a6abefe1b4b916ca51c3e958e40dc78c3661313e0ed2e77d, 224'h6404d8a332a837f2ab6bd13e3ee4aad1e9307d449e7f9b7d6332030c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{276, 1'b1, 512'h0392f8c2dc961605c5693d9452731b6a8292ff57d6995aeca0dad3117459668ec7809dc09cf154170fcd624be50000000026e3d92dfdf1a2abd09392468117c9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4eca73709a67c41603ca5af494c8132483ffc2e0bf171b52de5a5e81, 224'h2c79137cd2add3ce3a76792270e347221a3ad786eafc2682b39bcf95},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{279, 1'b1, 512'h81b675425e8c528a0a51b23413c8b796411a01b207e0bafc5bd2a46b05237be84abdae1ebd492fca053bf7e3133392720000000086ce63108f1dc5a3b34c575d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h49886a8c26c91d649cbfecda6ce8d1441e764c66f5d81dceedb6c5ba, 224'h4370d8bcd4f052fac9491d62850b6a6a85d5acc44d9248c3dff30bf2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{284, 1'b1, 512'h99f941e73ab790b224ce0a799133f6b04eb9bcfb2fd0ec84b8e7d5dca6ca50d2b1ae4d31c57e2e54f97f59b6a10d0758cfb3e46500000000909d4fabd9d1962a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3d243581c0874fd4eb4d80f896c5067429ad455314881951ab5ec6e3, 224'h0ec47aba08ccba88c1a6ddc289f595bda08dc2dd34d12dcefb68094d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{291, 1'b1, 512'he698cebca57a541614e179f28ba51cf82fa0fb4300f81df5fe22b635eb4441b496a36ad280999f503edded3ae1cab1700758b5ae80ce33dbf25c7300000000e9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h187fb026ade3ad16dd4b2813e8ebda433cb6cc3af1615bedf486a9e2, 224'h6fbee53fa884d296f34f7719f74919434d1b7090c485eeed2fb8fd6c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{295, 1'b1, 512'h391dffffffff5a981c0576acae266e7b35ecdfeddfeb6db903e9f4eab200dba039b146517f0c5b418d096addeab6d0962a6f77c2a2a552748b788c07796553e5, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5be0e0dfb26b1caa88f866504aa8e76f035a82abe00028d962bcfafa, 224'h3c3c1df06026123471bed324ca79c51b28b3d10b1ce877cef21b852d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{302, 1'b1, 512'h6e50953fea8dfead2fffffffff824e02147d010595358c98ec376055cb9ddc1dfe6d3874cf38e8a98ef0664fd3b10605bc14506eb7e46460c9db81b10e2f6730, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1caece75c8e31bb0c5cceb0842f23683b8557a97036574ea88ceeabd, 224'h645ad3276aaee22b693647f00dce5f91a03b678b789b667cd3b8e751},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{303, 1'b1, 512'h1539fd34220ed16ae0b8ffffffff88a04bebde47a3a94f1b86bc687c2ce7648caa7d42ac8693b5704e401b7c9f4864bbafe3bcf761d862739eaee02516a0d707, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3a7d582068aaecaba945203bc445b3312e5cb40886522987aced68d0, 224'h39b3c612b6743a13bb2ffb83514d690cfcb9a7055e3a993cb0863938},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{305, 1'b1, 512'hc3b630a45b21b937bf78ef4affffffffad33da42317364a1090ed4446da7738caefc807ed99c92f85a6f6ba946f99284d4b9793896bc5e0b6f93cf1b09b35a6d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h79cf893f66f7faa5ca08553ea03456107e7bb391a5e51260cedaea84, 224'h32e8e3509468da7216c59975d4f3d5493848a03f864b2332044e68d1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{308, 1'b1, 512'hcd86d593a60faa34608d5bcdb2e878fffffffff06003c116f812eecd35fc6f3cccc1dee24c5cb89cfe9d41b0defa4e5d16b1d9aa4897e6efc838a8a6dd5f22aa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h258dce916ef78b9d8a87beaf6edd35bcccc08c5de488586e1b7b749a, 224'h4ff500db4d665c7062179c099b2985a814f99fbfa44a3a709024d589},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 512'ha6d55690f7fe8dc6a67ac00e5f136dab1f6855b53643ffffffff2585eedbf8e7c3db326f7fed8c48851376d7b1a34dfd79aa6837d19b05becbe8b8d122d1baf7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7ed658c30f4a0dcc894c39f9320f59a185509ffee45eac6023577c7c, 224'h47ac94a501806d5adffea9fcf3ccd8cf79f3cc47eca9fe38fc4886b4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{317, 1'b1, 512'hbf0fafaf135ee4e03b991ef87e6e9377150ae255e043de57ffffffff10002deb92f4bf4c1770933d3137b0165ebcf81c8c3387c21457e0fe0c39c7c7947837b9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h537ec369b3f0d891e166f6c74e5d73dd2c4822210c5fe5f978c34072, 224'h0b183c48b5f6e69245cb76e1e2c39663eedfb74ba9538739ac495ff5},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{325, 1'b1, 512'hefe7f8f35a94b65eb3a9299658db8b8256f29f2df969035fe5769c11e85c9b7bffffffff61e57fc3e05c9a1eaf760ce1b13dc6ddc5516048677e1fcd420a6427, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h66cda58a5a6ddb9476e36dbad5df542be88d7e447bdc3dfe1d9e8b2c, 224'h0d99d387486a964ebab4e29bad583e46a5a200391d1065768a4e35fd},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 512'hc5c3daa9bce3e7422af1de2fdc992b34f5c8ef3fd448b45f2426e1677feaa86aa3ffffffff6e9d87ba471035c9beb5d2c94f3bb0dfb4c48298a8615840c621a6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3200761902825bd353908accd2be6b482645646971f96dc490706a37, 224'h3ed77899efdbe418370fa7998df3b7c924bed6864535277f805c894f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{330, 1'b1, 512'h3be3c1c0f8b8f6b9c476455ceee9edbf99283f1eab4a28ace9494eae8da166e4aa1d5def8affffffff3d69a06db8c19c0984bdd10df6ede19e4214183d3b0762, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h331a1a553494f8524adb4e8a722d558965fb703ae432bf3cbdb255c2, 224'h5ab6e3dee6a2516fc4e0ac88e6dfc81d2bc37c98949cc03e521d389d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{339, 1'b1, 512'h0477828c9cc5710ded82ab21dfa5887f29edfb47548a5a99ff8315da76be5f67922c0a5de1cb7448a3a79b214889ffffffff7dc823ffb5d2fbcda33e63489df0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h54d6d44373f7dfc98455a22cd39a0b320fabc33215216b37365b5a16, 224'h29cc690f2467c02e07bc416ad47204975af8c5c3346973f2b03ded3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 512'h17dfd1c9bfab4afc7d5ac126157041f4c4ca4a04aaf17c45e47857c384fb415e4362041ec3e91609325b7e4c9fb1a3ffffffff9d3efaa9406e392a0dea1ea309, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2f5048c9ef9f30da7cb3fe4624552200f9e57a46d79db0484a0d9cf2, 224'h06dad3a4682725852869a1a459bec865661e1a38a9e546eeaac7cb84},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{343, 1'b1, 512'h6ea638f8043673b9b6a79ff39b5d311774de5f4d697e5251ede52feecabba85d705f25c58b7c2efc844ce598d1428d22e4b3ffffffffc75b0ecb7283d80278f0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h43ee11a7ab62e2125e765c2ce5d4f84704183539810512268d87f195, 224'h65897e54025777659ee802b39c6bfd5ccc5706a9d1b38f95c078abaf},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{347, 1'b1, 512'h51ae80a63d993770d8a5957111af53dabdf3abb9cf9908bc162ded716d3b3c5af2924c076e87c96249a4d7650253ff5112f8a2e7d2aaffffffff66e0e9175efa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0b7b5aab8364dd4b11001a0b986d5aa4fb61ee720237417a7f63722f, 224'h7f13b411e645e819fed1b925ebe807d9560b44d0ba1b75bd2fbd1294},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{348, 1'b1, 512'h100c883756f36d7c944d934c08932a99a1c2eb9892cc39a13a80b22aadc526ad755265f9ebbc8d0c1ccd31240299c71604332ff56592b7fffffffff1224308a3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h505b974f8ecf07b60ffdbd2b2df9324de92b39476eb763a4c25f126a, 224'h1c36ed1dee772c724205f717c383f49a87a5bc3caa0ef81360f9d800},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{351, 1'b1, 512'h8a5409853b325b917b8a2aa1eb394767bb07fa82af11357e777f7404e0955bc9bb9cc5a918475c52df4772a1207e3ee4f3e3d3c8e68e84e10477ffffffffd35f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h24916961dd0d168c2878ca4fd065b81311c03b7f23f8416f4a23b14b, 224'h1e37e3c03b2333b33bbb2ebe05b031042af19315adfdccdfc8d078ee},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{354, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6239877430e268f1a3ada2c90357247c6ca6687f49023bed0fb5b597, 224'h355c60c09f0dacb9d74b7ccde71806c50fda8750c6ecb7abba910ac7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{358, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h2f6983b6e9f8ef96c2d981f69be54b06591ed73fe40c8a546b936a79, 224'h71bf57726c26c811d7625a9d851951c1fffe236b0eb3b896bc4c98ef, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{360, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e8f90a717714f0158d9521f18c14ae8c83bf1eeba115c46cbdabb20b, 224'h66f50ac13461c02da02edfe4296a1f543dde7b4359f905e04193d3cf, 8'h03, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{361, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h723bc0c9b7ce6ea784ec075036cede90452c76576bd8fb5be4dc0fb1, 232'h00cf405820d92f48552b551c7b11f49406dc892fd659971ae7f9e74b59, 8'h03, 8'h03},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{362, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00a0dcce127084f955a4e49a7c86b9b91b05ae7afd6eb07225a6541d88, 232'h00f10a1d4fef93934967bb6c5d8792bbd47ab3abb406899a00b1c91b4a, 8'h03, 8'h04},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{366, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h0091a85b3c5e90b409f6b8d3bca9117a54a40f4162b388bb9367fd6439, 232'h00f1cedf20ab52eb7154b7ea1f2934a9c8292906e18a0e572002cd2f7c, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=56b(7B), s=224b(28B)
  '{367, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00d1ca7a5c1aa086b2951c1ac14e005f0072fb28383973a05117f9652c, 232'h00ce523c05ebe94991c47fecd241d0a07e86c88ab3c620eae792aba3d1, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{371, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c2ae0e357a43f97549a725ae3704449051c96bf3633355c35b6eb7e9, 224'h6a84dfb6d4517d1de46b18786a506178724bf4ae4f9e418c75ab17ef, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{372, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c2ae0e357a43f97549a725ae3704449051c96bf3633355c35b6eb7e9, 224'h6a84dfb6d4517d1de46b18786a506178724bf4ae4f9e418c75ab17ef, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{373, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00961617d9855f202fd600b584abe94a46674927cfdc6333c5be56ce7b, 232'h0089b4150d9ccdfbd77e7682ca862c0c3e96d89c918b7d3b7bbb92ff43, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{374, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h008db53fe4168df43ee538bc9d758b8c26fa433fb0101bcbad039585de, 224'h2310dfc20835379ea406993036fd4bb0f67d14760e1eb414c32dd1f3, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{375, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h0b7fa61983e7a227f738847d457f3e8cf0a4085c312fb6dcec822570, 232'h00ee7434ce2ff3fbcc1d0960379876e9dd5bed28aad576eea233a44b0d, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{376, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h55b212919cd6886b13cd7a2556430ce442e86942f1bf6e4618ae363e, 224'h795c664ae960ee1106308b7dba91240ab0c3ef8beb7d0a4d7a102a7f, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b0},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{378, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h0c8e2cb5f6a903e1cccf3ac2d465f1d0dc3452237fd9e8a4df5d5341, 232'h00d044ca8ceecb54a1b951270971e5ab4eb226116c48c553499d1a4899, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{381, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00f49278419e4f506889b0168b1fce1f87ee5b61efa0e73c7833eeb29c, 232'h00b1b334f81be8f05f3b2e98d38b030cff57947b96135ec4465c5e53f3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h4e158ef86cc53054f1635c74e65508206048929315e097a59f1519e2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{383, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00f554014cc14f319c18f5fa6cd739249075ff35ba3b2afdab5329ef0f, 232'h00d2c501f25a704addbd85c0e022748956e5998d99c387fbfd343c89e0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c5221f3c2de0c6fbc07ff04150679b57f57512b814f413aebafe731},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{384, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00bcfa8db704aca56feb23bd4b4049213233aa652045a0a81a2e0da64c, 224'h091b359f7be7ae00a0e9777d9510f847430b5dfda878e66d4fb0d62f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h221f3c2de0c6fbc07ff041506dc71b5a312063d87beb4c30c289210f},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{385, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h009fd4d828ae98056be58fa69eaf9cde98ca0ed9b415d6463fa1864d9f, 232'h00b2a5e41f10e8789450217daafd259f204aed87b0e26100f43f7c5bad, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h443e785bc18df780ffe082a0db8e36b46240c7b0f7d698618512421e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{388, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e012c23c6867e9553313d0179e9db953de7c368cdb59abe05f1c52ba, 232'h00d352a57bb59c45159352c114eeb696ec3b79caa835ef5c2ae71ddcfa, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3ead55015c579ed137c58236bb70b0a2324e79109e2ffc964262f12f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{391, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h08842f19b114d16be27bb4b6971377ed6b1d0915e133a9ebf01674ee, 224'h4c97738b6912ff71553c4a747c782eddd9d2a20fbeae38864d217859, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{393, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h008fbe39e75bc4fd8a15e4b52e4bbebe2047d54385a7117e17a4d0b2b2, 224'h07abdb40824538e5787c718d6548583f523f6b5bbfa239a7f622c8a0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{395, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00816fdcf370827e3f7771564e1aa73ed73e62556deadad89711cef663, 232'h00edcda0ea42235f4c9a8c13f787351ffe5ceb32f15fc0ccb24e0a409c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{397, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h288f38fd77dd1603ff0275cb11cba280ae3408affa6a760f396f1a1e, 232'h00c84ca6fd772c6ac6cc523cc72c2e7e95eb6a36a66b5cca5a58ba078a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{399, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h75f007c11b93e6f46e9a815cb765990a8305d3ad8d22c76fe6b257cc, 224'h71b5c1951b5d464c66df7c290cf0a4f156bbf52f1e41a79dc63abce5, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{400, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h1255fb94a0f20e6faa2505c394cc3c39f07def4107127dffc4dacb6e, 232'h00ea73c1044544a1496560bd1b049ff615e68ae0d483220327569884e1, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{404, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e5462d3a838d4a14de96a7b0b1071eb622ae6e71ede8f95ff01c2121, 224'h368e3a90d8584e194616d3211a7541f6a0960339cab28e8bfd6b1dfd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{405, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h5d97670c1f121f7f1ba541505609f20143b312a7bb49d376690e1831, 232'h00c1b4567141a7b534e21bd2f706ae034169ab9c3f8536147904de8c5f, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{407, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h5a5cd1162388348734dae20e2235ae2c464adef0a196f9aaf02482ca, 224'h2ae94e8b9a024375036429b632ab485e02c5a9665b289b8a47bade8f, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{409, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00cf46960060453e55577f1bee6a9c4709e7cdcba45ca8020bb3536931, 232'h00ea4ec33309213864a1318aee0a86d8b6f0c1b9741cd6bd5dea4f4066, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{410, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h62f4eaf3797bdc3d5d8cfaa07b5af7060e131b183ca4eded4819e561, 232'h00bff3eadd7b55db2dc01bd20569e6c47c9212f9b2d6793795b51e4f6c, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{417, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b0, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{419, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b0, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{429, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h791624e5f234b8950d509d0b456ef6fa778b19dccd609d496b62a211, 224'h6c51e846fa53d03d42f798e6bb90954f9a48c1794b47e84ac97b460a},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{431, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h224a38e733ebd3fac274ecc50ecef2e7c3189be2b9d093a8dcc6fa3a, 224'h134fa5a4f923d296b3c6dd4683d249ccf0ad272890e4149c9a0d7415},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{433, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h689fce4b33d8212a663640a1ae0efaa7a7d7711beba719374fe634ee, 224'h04bd9981fa52293063076f0fd70fc31875d580ef94f020d2f95440e0},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{434, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h2a4287e01510e7fb5fed2e1ccc3f2a6929cf7d03850e49d7ae8a504a, 224'h355c3915f3fa9637dc8001438a8c04e15d14934cabd430feb0cb5ba5},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{437, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h54e6add8ac910e52c6228fe3980d8f586218334d8d859ba9a3329917, 224'h5836cc79ec88519eab4a6b2614c501628c9fee32fbafd93e32158409},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{438, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h1230d5409f379584b4d548b7bccba64baf81d512a9f2e6398c4e3a66, 224'h1937a298f8cbdfa85b8e6fcf0a12be4966d80270cade85a0c37ee6f3},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{453, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h5797c21c0162e42f69693c6c0244dfdf9218c01e9235760177b61a54, 224'h5452c887b27fb342a8a00d27579c7195dddb73df399233ed0dea567b}  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224R1_SHA512_SV
