`ifndef WYCHERPROOF_SECP224R1_SHA224_SV
`define WYCHERPROOF_SECP224R1_SHA224_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp224r1_sha224;

localparam int TEST_VECTORS_SECP224R1_SHA224_NUM = 224;

ecdsa_vector_secp224r1_sha224 test_vectors_secp224r1_sha224 [] = '{
  '{1, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'h2840bf24f6f66be287066b7cbf38788e1b7770b18fd1aa6a26d7c6dc},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{2, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'hd7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{3, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{93, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a0000, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=240b(30B), s=232b(29B)
  '{94, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 248'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb358463610000},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=248b(31B)
  '{98, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a0500, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=240b(30B), s=232b(29B)
  '{99, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 248'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb358463610500},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=248b(31B)
  '{114, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 0, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=0b(0B), s=232b(29B)
  '{115, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 0},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=0b(0B)
  '{118, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h72049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{119, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h02d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{120, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a488a, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{121, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb358463e1},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{122, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a48, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=216b(27B), s=232b(29B)
  '{123, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'h049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=216b(27B), s=232b(29B)
  '{124, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb358463},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{125, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{126, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 240'hff00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=240b(30B)
  '{129, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{130, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{131, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0170049af31f8348673d56cece2b26fc2a84bbe2e2a2e84aeced767247, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{132, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff70049af31f8348673d56cece2b28cee4c34a02667b2df86234be1dcd, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{133, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h8ffb650ce07cb798c2a93131d4d81a785bfd0d5b70f4de586ee5b7f6, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{134, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ffb650ce07cb798c2a93131d4d7311b3cb5fd9984d2079dcb41e233, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{135, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hfe8ffb650ce07cb798c2a93131d4d903d57b441d1d5d17b51312898db9, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{136, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0170049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{137, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ffb650ce07cb798c2a93131d4d81a785bfd0d5b70f4de586ee5b7f6, 232'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{138, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h01d7bf40db0909941d78f9948340c5b4b7a5fa6fca97e8a82091e08d9e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{139, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'hd7bf40db0909941d78f9948340c78771e4888f4e702e5595d9283924},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{140, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'hff2840bf24f6f66be287066b7cbf3961eb3abe80737bf48124ca7b9c9f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{141, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'hfe2840bf24f6f66be287066b7cbf3a4b485a059035681757df6e1f7262},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{142, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 232'h01d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{143, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'h2840bf24f6f66be287066b7cbf3961eb3abe80737bf48124ca7b9c9f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{144, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{148, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{149, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{150, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{151, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{154, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{158, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{159, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{160, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{161, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{164, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{168, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{169, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{170, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{171, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{174, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{175, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{176, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{177, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{178, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{179, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{180, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{181, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{184, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{185, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{186, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{187, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{188, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{189, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{190, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{191, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{194, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{195, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{196, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{197, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{198, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{199, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{200, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{201, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{204, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{205, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{206, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{207, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{208, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{209, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{210, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{211, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{214, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{215, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{216, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{217, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{218, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{219, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{220, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{221, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{230, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 224'h3116e1a38e4ab2008eca032fb2d185e5c21a232eaf4507ae56177fd2},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{231, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ce2afe20b684576fdd91b4b34168c9c011996af5b0eb85fa929f381, 224'h662af5ca651bffbc623c3a3b372779bd09e1948cd19188f5339a979d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{232, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00da573cf73aed174710c232155735248f8ebef696374647527da52258, 232'h00b251856b66a83c32bf0b7b81a01f1db4507e622125f301bd832a5ccc},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{233, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c368da86582b2c82b696b2f7c79027968f3fd25cbba9688cdc67b17a, 232'h00aba8e3c2ff1af9bb9c66ca88a3825a19ce17206e7a658ff47025891e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{234, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffcefcb57190d0b87efb789fb53407fd2c65c5ae3551da3eccf8ddd5, 224'h05c89b41238f1e1def8fbe8d4afebf20be077e82972f91297487e118},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{235, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2b98c67ebf6597b08bc7f1b73ff8662cf125e9700ec973ece9c6ff48, 224'h2e3f72a8f76e12c8cdf4487e0956c1ef4578e1da4d29d8db824d415b},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{236, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5794d70440f166904d24d0b910cd127c63a9eddca45a4d9032db47e8, 232'h008ba5d290834d9a0963122d928da902f7b03467396072180bb1801b43},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{237, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c29c70b0b21782d1c727f4907aef5641b6d6c6e7b2a1ebfa57794223, 232'h00aac2d3a02592f298dd3198e388425ec7a91d7e6be48248a64773614c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{238, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5c3ef3778c811e69ef0b0e370e45ec0d7eb88505c3e8ffb8c50b9993, 232'h00e06b5c6e47dc4da9e64fd21bc3e1da13cf7c264fa64ccb89da87387c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{239, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ed8f586563232cf15ebd014bd4f99727e337cfe4ce48694fe6748ec2, 232'h00fff779a3eca9513522908e252a2b4aab2060608e6cd2d4f1b8c696cd},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{240, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h64c084f6b775bbf7915c1964a68b0259629328598f13557872867830, 224'h2a6f3b289d130ec3d99e4caaf601497895a069c1a5a75b559ad28444},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{241, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2b514e9b0e0eb68adc01915abbee9fa21f3034be5581dedaa6b15982, 232'h00b8f71c5fdc68d698716bfc623b278216c0fcc0298497fc9c03db44e9},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{242, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e4103f4a8a814485b6b406fe8dd72206bad6a50e7126bc655c3d2285, 232'h009bcb99693284cac26e6641a861dbec24f9cc5dd7bb535339d09ac984},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{243, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009edfb833446ec8b6fc84eea34ee40a85b732e5c99da8abc8bafcc515, 224'h5052b40f9d407ae90003299cabe3e1a587b0558127cafb31de6b2638},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{244, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ad2647c8ff377798a6aeaed436d30c7b25fb52428829ce6424dd34e8, 224'h28f58671d77c86da302418c51e5ab86d137ba6ef4389722bc79b8751},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{245, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5dfc6fad385bdb24b2b70a64fd4253405c0028bb36f4793aa3bd31fe, 224'h1c210b74924171378992b03bb1bd78c5cfcfc879d2e5c736d35516c3},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{246, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h766bef46229695e6829dd12cd558369ec34519ba4a72dcaf6f73f7b0, 232'h00fc015ccdd1e943b910101607d81ff1398ca6a4d70c25832b02b221e4},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{247, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h120055f90ad1290c4c5fc5faf69b215139182c770d2b55e95712442f, 224'h01ac47f7446543d4003b039d9f54daa9d0799f98291a32df4fcd472a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{248, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f480591f6f40a25b37a035fd91954145ec342e593d09e142f25da408, 224'h5c6ba44ff52f52c51490743d9b650916be58d06d7c1fd99dfa2eab58},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{249, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h57daddb0cb6af939b1ea1aaf4bc72e56150c0c46a581827193e65d17, 224'h3bc37bde4e60b789ba86a054d37f1191e0814926c1a0100168d16c17},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{250, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3a74102bd1fc617018efc4fbc042e719a81b55830aac1f1dcdedec65, 224'h4bb9fe90015a45f31c8c95dda24f54fcdb64682c13f68d4da3d1abe0},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{251, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e3b6bb1b5beed048e0177e3e310fa14eb923a1e3274c0946f9275454, 232'h00e044e0494ff46573c37007e3efa3233588f1d103ced1823c7e87e7c8},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{252, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3c212b5a7e65d9af44643bd62fa42a9b9cffe6bdb623e9b9e4337156, 224'h29c8121a12427a324e5d551ff5a83d3c252e32257af2800d080817d2},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{253, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1630554989fffd0e35f2d9105623d73a543634c48000484c422272ca, 224'h214da487d5e51f73814dff80a08c77bd8a83a9889a1b26a5578ba954},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{254, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0a4609242f2193b94bc54f49bcf532a576e035cec50e043668574bef, 232'h00aa68bd67624d8812002bbb3a5f530594451372d4ab36896a2929c3df},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{255, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ef9ff446e8eef3e948f4129fe8804f81f5b7f116a5383f9e8bc359e4, 232'h00f4c7055bd98f4a7ea49d9574160eac167809f6a78b9dd220958dd0f3},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{256, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1a6c59d85d5b3120b28c0d30bc058a92dc725d8ef450c198cc3ca522, 232'h008b17fefc8ab1ff0bb37a93446453d40f65bc2cb9636b11207f5c90a1},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{257, 1'b1, 0, 232'h008bf7e792f7c86877f1fd0552e42d80653b59e3a29e762a22810daac7, 232'h00eec615bbad04b58dc2a7956090b8040bb5055325bba0aa8b3a5caa6f, 120'h00e95c1f470fc1ec22d6baa3a3d5c1, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=120b(15B), s=232b(29B)
  '{258, 1'b0, 0, 232'h008bf7e792f7c86877f1fd0552e42d80653b59e3a29e762a22810daac7, 232'h00eec615bbad04b58dc2a7956090b8040bb5055325bba0aa8b3a5caa6f, 232'h00fffffffffffffffffffffffffffffffefffffffffffffffffffffffe, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{259, 1'b1, 0, 224'h2646ff36d9697aaaed0d641117f94f60e138bab8e9912b558ae0a818, 232'h00ca48e45a33550c1b5bd20a00e4d9df3033c03222e87bd96a8197f2dd, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3b},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{260, 1'b1, 0, 232'h00ea3ea2873b6fc099bfd779b0a2c23c2c4354e2fec4536f3b8e420988, 232'h00f97e1c7646b4eb3de616752f415ab3a6f696d1d674fb4b6732252382, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{261, 1'b1, 0, 232'h0092ae54e38b4e9c6ae9943193747c4c8acc6c96f422515288e9698a13, 232'h00e8f3a759a1a8273c53f4b4b18bfcf78d9bb988adb3b005002dbe434c, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 232'h00bf19ab4d3ebf5a1a49d765909308daa88c2b7be3969db552ea30562b},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{262, 1'b1, 0, 232'h00b157315cc1aaeae64eb5b38452884195fdfe8a15fb5618284f48afe5, 232'h00e1fbbaad729477a45f3752b7f72ad2f9cd7dce4158a8e21b8127e8a7, 8'h03, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{263, 1'b1, 0, 232'h0087d9d964044b5b16801f32de9f3f9066194e8bf80affa3cb0d4ddb1d, 232'h00b5eb9b6594e6d1bcacd0fd9d67c408f789dfb95feb79a6e2fb9c4cee, 8'h03, 8'h03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{264, 1'b1, 0, 224'h461b435af09ede35e74dac21f9af7b1b9998213039f8785d4a4905f5, 224'h18b89bde69de34a482638461d09386e7193ca90ca5b3038e2a3885d1, 8'h03, 8'h04},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{265, 1'b0, 0, 224'h461b435af09ede35e74dac21f9af7b1b9998213039f8785d4a4905f5, 224'h18b89bde69de34a482638461d09386e7193ca90ca5b3038e2a3885d1, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a40, 8'h04},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{266, 1'b0, 0, 232'h008093af8db04b3dd2e7c3c59bb64a832c2fb8e8e141bae7ba1534950a, 224'h10c5e87aecbd1fcdfc36cd18d41b3238b2ac613eb7c9de988d881816, 8'h03, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c6f00c4},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{267, 1'b1, 0, 232'h00c6d71f4ba0933f1269f7d6df83fd0c9c67254f101dcc126dc15faa3e, 224'h3c45dc9fedc71c9f2b0dd1b12b656241f5e335066f3f925bdbcfe98f, 16'h0100, 232'h00c993264c993264c993264c99326411d2e55b3214a8d67528812a55ab},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{268, 1'b1, 0, 232'h00beb9d8dcba48146b9032688ecea947a231e7d0e6ce17d76b56ed6348, 224'h35503f3b4af414870ef03383784b1d846b3e07b8e9fc2d6190a3bfda, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{269, 1'b1, 0, 224'h1955ba3f90e7a739471a5d182b594c9747eb49d5356203f3bb8b939c, 232'h00807d88ce3a0885bfa5b5b7f6e9beb18285e7130524b6c1498b3269ee, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{270, 1'b1, 0, 224'h5cb9e5a5071f2b37aa3a5e5f389f54f996b0bc8a132ecb6885318fbf, 224'h4ec5f8b93d8bf2a3b64fa7cac316392562c46567963c43a69f7a37fd, 16'h0100, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{271, 1'b1, 0, 224'h7b34ef8723a4309c0fa8a7ec3a783477652a82892370f6763314fe7b, 232'h00dee663853071e35fd3c76f991d7843c5e168ca659b93bd6015518fba, 104'h062522bbd3ecbe7c39e93e7c24, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=104b(13B), s=232b(29B)
  '{272, 1'b1, 0, 224'h03f26a9c13979cf5d090ea25dc966398022ceec31504abc4b10f7676, 224'h7d577dcf47e10e384c6b9a229a455a9fd33e54fe7960b8b0160aef16, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c29bd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{273, 1'b1, 0, 232'h00b671296dd5f690502e4b1500e4acb4c82d3aa8dfbc5868a643f86a3c, 232'h00a46ba8c3a7b823259522291e2416232276cca8503cc8dbf941f1d93d, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{274, 1'b0, 0, 232'h00b671296dd5f690502e4b1500e4acb4c82d3aa8dfbc5868a643f86a3c, 232'h00a46ba8c3a7b823259522291e2416232276cca8503cc8dbf941f1d93d, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{275, 1'b0, 0, 224'h76e34b57a8c61df59cb0b7921cec6e5422344033f7accb7b3179e682, 232'h00cefd0a848309d1decf98a3b9e333691b95c17821cb681137630c02e2, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{276, 1'b1, 0, 224'h51839e545c872f4a381f278ed5b4c24cf38aac77b02953405618bf27, 224'h394e41226594c499db6a7dd7a6901bda5e6474b1ffa10a6567210010, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{277, 1'b1, 0, 232'h00a3ec90053d1e100815d1becfe96c9b3646e52df794f6b03b766a7574, 232'h00c3b7e17e73acc8cefe71b6eb13d4f1c94c57e58bee43c69d9d41a964, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{278, 1'b1, 0, 232'h00b5c09b4851a67371eee7bbf02451e5208c40de61bc1a33df2710b384, 232'h00dcce4e5b83c32a800e8de28fa936d582cdcad185e894caac797f1d14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{279, 1'b1, 0, 232'h00941e283be31300bfd4f6a12b876fd3267352551cc49e9eef73f76538, 232'h00c115e5fe3b92f643c6cef1c58f3f8657574d1f64957d4880995cde83, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h008ac44bff876cbf7e2842eec13b63fcb3d6e7360aca5698f3ef0f1811},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{280, 1'b1, 0, 224'h43c9ccd08a80bca18022722b0bdcd790d82a3ef8b65c3f34204bb472, 232'h009ee1c1f00598130b2313a3e38a3798d03dac665cff20f36ce8a2024a, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{281, 1'b1, 0, 232'h00d958e418fad1c5ea5c923e6185e03ed5539d3f5f58dfac8bb9f10459, 224'h6997e408c97be5fdc037a5c004389d4b97eb1f54635e985853c1f082, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaa0f17407b4ad40d3e1b8392e81c29},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{282, 1'b1, 0, 232'h00d629b434c9b5d157bd72e114fd839553f7f0e94600934a0a49e59aa4, 224'h713a13c01775e75e2ebae75d9e29d2506184177b7dd0868693873596, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d1be91557d866ad5f2945b14ec3317bc43c1338fd06af6496201cce2},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{283, 1'b1, 0, 224'h3d2e9bb9a712bf3ad42ac30659fdbda9be9956537f9f37cd05f0ff37, 224'h7d5982d6d9266d774942c44d9eb3501051d3b9688610131e7856ef36, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7ac54a381d9bd3f2698359d6f658b5e4167d15a75b576e82d2efbd37},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{284, 1'b1, 0, 232'h00a0be2f10144b9b42b016f1bd9fca30e4c24aae4775596c7cdb07ae60, 232'h00d60ff3a70f1541631f6087d3f3b3fe376d2305b50b94821106412479, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h4fbb063e82402e16fe14edda4d7986b0b88344a1f53b0e2684ee7e31},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{285, 1'b1, 0, 224'h4d74397a586c8ac5e326bed03720bde7037e4a07aee7209f70493cab, 224'h106778bfd081d17ab6dcb8fd8a454962941c26ecc19cda9fb77719db, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d3be5f50d726f99b8ac44bff876bfe78dd7ae630d227ef0ba87ae39b},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{286, 1'b1, 0, 232'h008c2f149b1738243f81a6f12135395a2ba2718863622e66e33efc241f, 224'h5638cf6ae9cfb39578cf3a719702052e5e9e940216c5136dcb6ef085, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00e5f50d726f99b8ac44bff876cbf710e47f9087d1afdfb1dab6d6daf1},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{287, 1'b1, 0, 232'h00ad5227e48afaa165e7b97ef8210687556e10643fda8a377aaf4f5bf4, 224'h12e86d4ae55f4460aba6a932f307ee78efdc136e9a3df6313100bf4f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00cbea1ae4df337158897ff0ed97ef0b261e681f654be23a7011518ba5},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{288, 1'b1, 0, 224'h3fb94a3165ecdef43fa27907ed075caf52c25420ac7bc7bb90408992, 224'h023c4d7b4775b591ae223dd4da9ceaabd73b9743ddab8b40576e393f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d726f99b8ac44bff876cbf7e28422aa07ec3cb1d9472bd704f4029f0},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{289, 1'b1, 0, 232'h00e45fcf0a7f4dc2a308dc7868251423fbf71a205a9546850a01a732fc, 232'h009a73ca4d41175076f2f362b276ecb0ccdb6e0bb30c4a1b35c2e3ed82, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h009720b755413cca9506b5d27589e58ac4bed856762ba7ae20ab5b43cc},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{290, 1'b1, 0, 224'h3c59e13982fd9c1a45991b1e9d79e939a52a62ca479764f1477e2813, 224'h1b004c9bffd7f00c05e3168c625cc93ab7a0f1ba8d6fa26a4d5162cb, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2e416eaa8279952a0d6ba4eb13cbfee69cf7bcae437232fbfa5a5d5b},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{291, 1'b1, 0, 232'h00c6b8ff152d7a1b7a99ce3483bdeaaf5bd2ce64dc6b0f89cf3544b87c, 224'h053ab6cf9cb510dc1440ab4e412a167f4c69365fcfc97f31d5ba4581, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00c56225ffc3b65fbf142177609db189ab5bd013246f19e11ca5b5a127},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{292, 1'b1, 0, 224'h7c0772fb6553c0ec0dd1f73b5db380764d9f2f7afb4eac1e774dacd5, 224'h6e2e5de0db63bf03cf9675eae6d2dfe5424e79ab394951c9b60ad5df, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00a7dd831f4120170b7f0a76ed26bc4ea9cc9e1a70048c1bb5f0a55437},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{293, 1'b1, 0, 224'h4108e0ccd47cba09fb7ed4d9f3455823780965157861c1bf8f93d34b, 224'h46d6fdb71e9e89adaae71376b13fd17644b11eed00d498783da0ba1a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{294, 1'b1, 0, 224'h2f2da40a1b72f67ba63613a243119c41c7252839cf106e86b5d8e6e3, 224'h5a1e0e2fc49b4f316f0c0e7236785749eb34ce923c23aef330af8733, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00855f5b2dc8e46ec428a593f73219cf65dae793e8346e30cc3701309c},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{295, 1'b1, 0, 224'h7dc09710f4f586af05b08f0c9dcd48b1308733c97767fc286d1c7283, 224'h4353a704c7950b8f4a11394bc8db06adccf19d8ed95c7f214a173137, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{296, 1'b1, 0, 232'h00dbb439e2c3e9d1822b94ccc7d98c9fcb668e65dd6a759ad2dfdcd328, 232'h0082663234e6da512d7d7d5fe79156ad0e19ffc62d618e3cf48276106d, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0084a6c7513e5f48c07fffffffffff8713f3cba1293e4f3e95597fe6bd},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{297, 1'b1, 0, 232'h00e012dc20cca5bd2adfaa27f57419596ce09ed0f18a9148e30a0f6ed2, 224'h55beca1b5e3e2485ef9537ae48a67b72dbcf6d7b33372023a5c443e8, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{298, 1'b1, 0, 232'h00c510ab34abd4855c54d62407abe6ca090c73ba49aca9de9bf117bca2, 224'h42b3b00c272c22681af7c255120fac148ad73c81b47846e4ad2f5627, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d8ea27cbe9180fffffffffffffff3a43fa3662a899627950d4eb64bc},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{299, 1'b1, 0, 224'h08a6e167536a47aaa224fec21ce077642efdb97d93ae16b9672279f4, 224'h33fb9f1abb25f2c0c3e6008ac857ede4a89ca8d9d08b8996614969ac, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{300, 1'b1, 0, 224'h1a83e185fcf30e6c69cf292e497d63cc04e6fd07cb9365a74be3c39c, 224'h6b2d56247df49cf94176c4e8efc84ec710cd0d614dd066c16f6ad3e0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00bfffffffffffffffffffffffffff3d87bb44c833bb384d0f224ccdde},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{301, 1'b1, 0, 224'h2d59efd841a44b83fd42e6a2984a53fa93ad242c11678f92202cccfb, 232'h0095bcaf0b2f6eb0e6d4d83e3260e037d3dc0e48ab6c4141ce6b56cad0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{302, 1'b1, 0, 224'h1161c7add6f67f995b93e19eb18bd5e73fd71d6bb10dceef0b792e9c, 224'h08c44cef9826b4ed67508c09d07ec857a0ea49ed1a7f1fa2c74cb838, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{303, 1'b1, 0, 232'h0084dc3d2ebfcf3480713baeff30ad0781bc8c4d06ab6ddd4f7f1045af, 224'h7570537c5d71a78b1a041aca0fe35f642824abda8c3ff2e9fcf5c8cb, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0096dafb0d7540b93b5790327082635cd8895e1e799d5d19f92b594056},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{304, 1'b1, 0, 224'h1767574e645c550ef3d353f76d4428f9616ac288b36378857de33262, 232'h009fe09825a57f3a0ec11189f4560272297ab6d5e095401febb60d0dc9, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h1ef359e4bd146f63d8155c5c2523fa3353c9820f84f28150bad3819a},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{305, 1'b0, 0, 224'h1767574e645c550ef3d353f76d4428f9616ac288b36378857de33262, 224'h601f67da5a80c5f13eee760ba9fd8dd585492a1f6abfe01449f2f238, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h1ef359e4bd146f63d8155c5c2523fa3353c9820f84f28150bad3819a},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{306, 1'b0, 0, 232'h00e2ef8c8ccb58eba287d9279b349e7652cca3e7cda188a5f179d77142, 232'h00f87594f3664c0faf7b59670e353a370d1d68ad89d6a1e246b4d03bee, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{307, 1'b1, 0, 232'h00b8bf3ef9646abfffb84220104ec996a92cef33f9328ec4cb1ea69948, 224'h4fea51a0de9e9d801babd42ca0924b36498bc5900fbeb9cbd5ad9c1a, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{308, 1'b1, 0, 224'h286e80429c8796dcd885d95f960d209fed19f87e2ce423d166c8e220, 224'h2e30882c09970d5dd58b67e5bb80affec74248a9cb4a783384c8b6a0, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{309, 1'b1, 0, 224'h5599a3faf96aba7302bd3d98cfde69525b7292762383f4a0b5c31039, 224'h3faa45feb6c35d2b7bf25ffc633c420ebfc4e715765302c5a11ac793, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{310, 1'b1, 0, 224'h5b5234b8db6bbd396eae7d1ca4e6d877824c98cde9fbfab34b6b8ccb, 224'h1f38ae9f87adc3e6d2474eb5e3cd9aeff0927320214be550f5e62ed4, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{311, 1'b1, 0, 232'h00aced4ea8949e5ae37ef2f5eb5e00675d08e17c34be6677b0f269b672, 224'h5e3ad0af49ebfff415ee4f2a838ead1f84cafaa652c17acc26130725, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{312, 1'b1, 0, 224'h3e8c1bcc16195e8769e25d4c859807dffe178bed5bca9db06efa1532, 224'h4e3b53b3048b8ccd8cdc1265be240c8ee204060486a99ad31eaad3a4, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{313, 1'b1, 0, 224'h24819323b7be8ab0910f7f33bd2f7669c44b13f09479965e95287d13, 232'h00b0592345beafbfdb8cf3629269bdd817728d5d5cd3c28bc6c6414a70, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{314, 1'b1, 0, 224'h44cf57bac30a83da39f90bf3faacd52211a70fb92547db7778ea6c81, 224'h2b3fd1bf14688d2770c50cd5a890a3807ba0e8612136a1b11e030f82, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{315, 1'b1, 0, 232'h00dc17f1001d326127f7375cffa70b7530bca4da1040dc43d0044aaca0, 224'h7a146f04c5294cfe7e1ed587da55bae70b7fa8e32f6aa800314d01dd, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{316, 1'b1, 0, 224'h68e2d7088eac18ba775bf68c5c509e86afd6f93451b4e4ee1d73e277, 232'h00e24ff4e27ef6c519db676d822c5db040482888013c8f3881bc9ac65a, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{317, 1'b1, 0, 232'h00cd4171adcb8be75e7734061a048b2bf228d167c2742d27f854392046, 232'h00865eb958ebd320ba87662ad3ac7af568c6be0f09be090bcfe083b3e5, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{318, 1'b1, 0, 232'h00eefdf99ab69d1888772cabe21d406045e1beab82761a7040beeb7ed3, 224'h59718c889af80f22f320fbe662d5ea0f65dfb4a5589c294ce5b73359, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{319, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{320, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 232'h008ac44bff876cbf7e2842eec13b63fcb3d6e7360aca5698f3ef0f1811, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{321, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{322, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 232'h008ac44bff876cbf7e2842eec13b63fcb3d6e7360aca5698f3ef0f1811, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{323, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h2770403d42b7b45e553308d1f6a480640b61cac0ae36665d6f14d34e, 232'h0085506b0404265ededf9a89fc7c9c7a55c16c5b0d781f774de8f46fa1},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{324, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00b68da722bbba7f6a58417bb5d0dd88f40316fc628b0edfcb0f02b062, 224'h5c742e330b6febadf9a12d58ba2a7199629457ef2e9e4cecd2f09f50},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{325, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h01ec1ff15c8a55d697a5424d674753f82f711593828368d2fbb41a17, 224'h20d9089db7baf46b8135e17e01645e732d22d5adb20e3772da740eee},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h3e46e9ba4dc089ff30fa8c0209c31b11ff49dbeec090f9f53c000c75, 224'h6f2e3b36369416602bca83206809ed898fcf158a56c25a5474143f68},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{327, 1'b1, 0, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h77b38da37079d27b837613ac3e8248d66eabd5d637076c8e62c7991e, 232'h00d40cd9f81efc52db4429c0c1af7c1d8a22b6c7babbe7fbd8b5b3f02f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{328, 1'b1, 0, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h008c03b32c166c0c8b99d7f876acd109447efb13f6b82945e78d51a269, 224'h657568f1a0a8bd7df5ffa43097ebb2b64435c8e3335bcaafc63f9ed5},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{329, 1'b1, 0, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h00d199a375253d30f1d2b4493542e9934f9f1f8b0680117679f5bc4ad2, 224'h11419ddbf02c8ad5f518f8dac33f86a85e777af51a034132e2767a6d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{330, 1'b1, 0, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h008ff82699e2e82870be9cfdd8a408bb34f8f38a83a4ac8370f18f2bc8, 224'h7e5008fab6a0d4159200077ef9918dad6592cd8359838852c636ac05},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{331, 1'b1, 0, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h3f3b60b529ae0f950c517264adf2e481616bc47416742d5103589660, 232'h00f731ebe98e58384b3a64b4696d4cc9619828ad51d7c39980749709a6},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{332, 1'b1, 0, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00dc11ffdc6b78754a335f168c4033916a2158d125a3f4fed9dc736661, 224'h6dd84364717d9f4b0790f2b282f9245ecb316874eac025600397f109},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{333, 1'b1, 0, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00a59b25b786d55f26b04dfe90ee02a6bde64ed6e431dc9fbdc3ab360e, 232'h00fc14b5ad20f39da9900e35437936c8626fccf6632e7a3d9e587e3311},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{334, 1'b1, 0, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h2eda1f96c1a6e3ad8a3321ce82cbb13a5b935b501abf6c06f7fd2b3f, 232'h00e81050c3e5f53a3c7b9d0bdb9ed92a326dfeac44791ba1abe4d6e973},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{335, 1'b1, 0, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h60f5e093fda08fc14ac99d820a18ad1370c58150bea0aca24fc6db9d, 232'h00c2220a0ebbf4896e68fdb5bd824f88291c1c862b916f9c4af87f8f5f},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{336, 1'b1, 0, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h2ead37846a5e36a490b75140bdc7b636c6e9f6d8f980f6fadb08f769, 232'h00e1fe130ae1798c196d7be62c7a5ddb3168cf4b8d48b6b6b4dc94ab3b},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{337, 1'b1, 0, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 232'h00a8a4c9416d72c860573d073281cb08c86ad65313f06b15a329e82eb2, 224'h5a6edd2f0816b7263d915d72c67d50a854e3abee5cde1b679a0cef09},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{338, 1'b1, 0, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h576bb86c517bfecdc930a4c8501725548d425afbb96d93f5c1e2a0e1, 224'h77248c5ecd620c431438c50e6bee6858091b54a87f8548ae35c21027},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{339, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h34e41cba628fd8787ba1a528f6015d2cae015c1c9a866e08a7133801, 232'h0083d422ffdd99cc3c6d7096ef927f0b11988d1824e6e93840ff666ccd},  // lens: hash=0b(0B), x=224b(28B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{340, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h2558a42e79689244bccd5e855f6a1e42b4ff726873f30b532b89ef53, 224'h07f9bd947785187175d848b6e2d79f7ab3bbc1087b42590b0cfb256a},  // lens: hash=0b(0B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{341, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00d5fe7dd5fb4fd1ea5ce66c0824f53f96ce47fd9b6c63b4d57827fd17, 232'h00bce5bc3af705afaacb81bfa6d552d6198962fece9fba41546c602ddc},  // lens: hash=0b(0B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{342, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 232'h008c1da2f07cdcbce4db8067b863468cfc728df52980229028689e57b6, 224'h32175c1390a4b2cab6359bab9f854957d4fd7976c9c6d920c871c051},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{343, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 232'h00e46d4f11b86b5a12f6fe781d1f934ef2b30e78f6f9cc86a9996e20c0, 232'h008351974b965526034a0ccef0e7d3bc13d91798151488c91533143f7b},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{344, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h305ccf0b5d0cf33dc745bb7c7964c233f6cfd8892a1c1ae9f50b2f3f, 224'h785f6e85f5e652587c6e15d0c45c427278cf65bb1429a57d8826ca39},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{345, 1'b1, 0, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h0e4fde0ac8d37536505f7b8bdc2d22c5c334b064ac5ed27bea9c179e, 232'h00c4d6bf829dd547000d6f70b9ad9e9c1503bebcf1d95c2608942ca19d},  // lens: hash=0b(0B), x=200b(25B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{346, 1'b1, 0, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00818afcaf491da9d08a7cc29318d5e85dce568dcca7018059f44e9b7e, 232'h00bf32a233d5fc6ed8e2d9270b1bdad4bbd2a0f2c293d289bd91ffbcf3},  // lens: hash=0b(0B), x=200b(25B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{347, 1'b1, 0, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h0e05ed675c673e5e70a4fdd5a47b114c5d542d4f6d7a367597d713ea, 224'h26d70d65c48430373363987810bdcc556e02718eab214403ae008db4},  // lens: hash=0b(0B), x=200b(25B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{348, 1'b1, 0, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00ab7a19eecf63e9668278963b65236b2768e57cae0e268cb86a0ddda1, 232'h008829f5d3a3394f9467ba62e66ef1768e3e54f93ed23ec962bc443c2e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{349, 1'b1, 0, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h17111a77cf79bead456ed86a7d8a935531440281eb8b15a885e341c0, 232'h00fdc3958d04f037b1d4bb2cee307b5201be062e0d4e089df1c1917668},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{350, 1'b1, 0, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00acafa1e33345eeba0c338c2204b4cd8ba21de7ec3e1213317038e968, 224'h0b42fbbaeda98a35da0de4c79546f3a0f7d9dec275d2cd671f93c874},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{351, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00a3fe71a2a56f554e98fd10a8098c2a543c98bc6b3602ef39f2412308, 224'h5d1d68f9a870ef2bc87484b3386549fae95811ab72bc0e3a514720da},  // lens: hash=0b(0B), x=232b(29B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{352, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h132f7625704756c13f2bfa449e60952f836f4904660b5b1da07e5a9f, 232'h0082b4abafc40e8fd19b0c967f02fff152737ce01153658df445c4d7b7},  // lens: hash=0b(0B), x=232b(29B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{353, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00f36a8347c6fe0397a1161a364cbc4bdfb4d8b7894cbaa6edc55a4ff7, 232'h009c9c90515da5e602d62e99f48eac414e913dd0b7cbf680c1a5399952},  // lens: hash=0b(0B), x=232b(29B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{354, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h2125ecc08e52e9e39e590117de2145bd879626cb87180e52e9d3ce03, 232'h008f7e838d0e8fb80005fe3c72fca1b7cc08ed321a34487896b0c90b04},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{355, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h00e485747ac2f3d045e010cdadab4fd5dbd5556c0008445fb73e07cd90, 232'h00e2133a7906aeac504852e09e6d057f29ab21368cfc4e2394be565e68},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{356, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h00a4de0d931ddab90e667ebc0ad800ce49e971c60543abdc46cefff926, 224'h550816170bd87593b9fb8ad5ed9ab4ddb12403ff6fe032252833bac4}  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
};
`endif
