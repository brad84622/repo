`ifndef WYCHERPROOF_SECP521R1_SHA512_SV
`define WYCHERPROOF_SECP521R1_SHA512_SV
typedef struct packed {
  int           tc_id;
  logic         valid;  // 1: expected pass; 0: expected fail (zero/oversized)
  logic [511:0]  hash;
  logic [527:0] x;
  logic [527:0] y;
  logic [527:0] r;
  logic [527:0] s;
} ecdsa_vector_secp521r1_sha512;

localparam int TEST_VECTORS_SECP521R1_SHA512_NUM = 316;

ecdsa_vector_secp521r1_sha512 test_vectors_secp521r1_sha512 [] = '{
  '{1, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h01d74a2f6d95be8d4cb64f02d16d6b785a1246b4ebd206dc596818bb953253245f5a27a24a1aae1e218fdccd8cd7d4990b666d4bf4902b84fdad123f941fe906d948},
  '{2, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{91, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf86450000, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},  // OUT_OF_RANGE r_len=67 s_len=65
  '{92, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'hb5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac10000},  // OUT_OF_RANGE r_len=65 s_len=67
  '{96, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf86450500, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},  // OUT_OF_RANGE r_len=67 s_len=65
  '{97, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'hb5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac10500},  // OUT_OF_RANGE r_len=65 s_len=67
  '{112, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},  // r=0
  '{113, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{116, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004c4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{117, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h002ab5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{118, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf86c5, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{119, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318a41},
  '{120, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf86, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{121, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00004223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{122, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h000028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318a},
  '{123, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0000b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{124, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'hff4e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{125, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'hff28b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{128, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},  // r=0
  '{129, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{130, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h024e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbe97b3367122fa4a20584c271233f3ec3b7f7b31b0faa4d340b92a6b0d5cd17ea4e, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{131, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'hfe4e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbf4d826580ab145752e852a6e91512b78178047879e9714a4ae1bc74298aaa7223c, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{132, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00b1bddc11bc17347621c4ecc6003d861a7d07d3854f08e4421bc241c8b538a00410d65320718f8af465fb099025b7cae2184402aea8df4f13a328c90648c42079bb, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{133, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01b1bddc11bc17347621c4ecc6003d861a7d07d3854f08e4421bc241c8b538a0040b27d9a7f54eba8ad17ad5916eaed487e87fb8786168eb5b51e438bd675558ddc4, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{134, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'hfdb1bddc11bc17347621c4ecc6003d861a7d07d3854f08e4421bc241c8b538a0041684cc98edd05b5dfa7b3d8edcc0c13c48084ce4f055b2cbf46d594f2a32e815b2, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{135, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h024e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{136, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'hfe4e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{137, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01b1bddc11bc17347621c4ecc6003d861a7d07d3854f08e4421bc241c8b538a00410d65320718f8af465fb099025b7cae2184402aea8df4f13a328c90648c42079bb, 528'h0028b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{138, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0228b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba09a7b6ac4ecd0410b4722ca75ba197a403a0a1f9ee0e7b391b0649fda1d3969eeca},
  '{139, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'hfe28b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a5d85db5e551e1de70233273282b66f49992b40b6fd47b0252edc06be016f926b8},
  '{140, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h00d74a2f6d95be8d4cb64f02d16d6b785a1246b4ebd206dc596818bb953253245f5fd61bc296eeee8b245d018b8edd8f659631962ad7a1e8b5fe56cfdd0157ce753f},
  '{141, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'hfdd74a2f6d95be8d4cb64f02d16d6b785a1246b4ebd206dc596818bb953253245f6584953b132fbef4b8dd358a45e685bfc5f5e0611f184c6e4f9b6025e2c6961136},
  '{142, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h0228b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{143, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'hfe28b5d0926a4172b349b0fd2e929487a5edb94b142df923a697e7446acdacdba0a029e43d69111174dba2fe747122709a69ce69d5285e174a01a93022fea8318ac1},
  '{144, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h004e4223ee43e8cb89de3b1339ffc279e582f82c7ab0f71bbde43dbe374ac75ffbef29acdf8e70750b9a04f66fda48351de7bbfd515720b0ec5cd736f9b73bdf8645, 528'h01d74a2f6d95be8d4cb64f02d16d6b785a1246b4ebd206dc596818bb953253245f5fd61bc296eeee8b245d018b8edd8f659631962ad7a1e8b5fe56cfdd0157ce753f},
  '{145, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // r=0, s=0
  '{146, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},  // r=0
  '{147, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},  // r=0
  '{148, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},  // r=0
  '{149, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},  // r=0
  '{150, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},  // r=0
  '{151, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},  // r=0
  '{152, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // r=0
  '{155, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{156, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{157, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{158, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},
  '{159, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},
  '{160, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},
  '{161, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},
  '{162, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},
  '{165, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{166, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{167, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{168, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},
  '{169, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},
  '{170, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},
  '{171, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},
  '{172, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},
  '{175, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{176, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{177, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{178, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},
  '{179, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},
  '{180, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},
  '{181, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},
  '{182, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},
  '{185, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{186, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{187, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{188, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},
  '{189, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},
  '{190, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},
  '{191, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},
  '{192, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},
  '{195, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{196, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{197, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{198, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},
  '{199, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},
  '{200, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},
  '{201, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},
  '{202, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},
  '{205, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{206, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{207, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{208, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},
  '{209, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},
  '{210, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},
  '{211, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},
  '{212, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},
  '{215, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{216, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{217, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{218, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386409},
  '{219, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386408},
  '{220, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a},
  '{221, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h01ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff},
  '{222, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},
  '{231, 1'b1, 512'h855fca3bb1b1130caf142425cc518a978f80236308b93cbe02d2455f14689f8393e55b9c35dc2b0388bce30b12742435c6b57aa7d5e63f2f2563325ea3bc9237, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00b4b10646a668c385e1c4da613eb6592c0976fc4df843fc446f20673be5ac18c7d8608a943f019d96216254b09de5f20f3159402ced88ef805a4154f780e093e044, 528'h0065cd4e7f2d8b752c35a62fc11a4ab745a91ca80698a226b41f156fb764b79f4d76548140eb94d2c477c0a9be3e1d4d1acbf9cf449701c10bd47c2e3698b3287934},
  '{232, 1'b1, 512'h0000000001b99889c891f2468c618149cb6865b933cca31eddb353de09746b540616ba69c5f5ff992c6d6177427daf1cb46a4c5c08625263a615fbf3eeaae178, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01209e6f7b6f2f764261766d4106c3e4a43ac615f645f3ef5c7139651e86e4a177f9c2ab68027afbc6784ccb78d05c258a8b9b18fb1c0f28be4d024da90738fbd374, 528'h01ade5d2cb6bf79d80583aeb11ac3254fc151fa363305508a0f121457d00911f8f5ef6d4ec27460d26f3b56f4447f434ff9abe6a91e5055e7fe7707345e562983d64},
  '{233, 1'b1, 512'h7800000000c52e48c315d5276f18d994c345b5805aa02872c29105d1bf75f152042a782853b4a3850822714434fefe3db00a19bc7eb84029869a7c1dca47ce71, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01c0832c973a455cac48a4439659aa21146036c52ec1514121c66714348a1c0e2c7099a2466d9acb49325a0cb509e5dff2efbcd90369d3027cbb7dca58a134278d05, 528'h00a426c063ab5cc6af20dd1ba8a519fac910183561598e67c0929e25f9c3aaeb245c5647fba21e30c103304dc6f49e6dec68a7833533e4e5448240bde023fe201eb9},
  '{234, 1'b1, 512'had9a00000000987c9531c475b0236659fdd3dd795473bafb8f0753bcaa4bea4e6418f79cba317764c48fdfd9461986dcf668f250be9ed2b7b75afaac70ccf0ec, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000d01cde64dda4dbcef1a9b924779598217b97eb688d9b4a4fd20d1b81ff0bb870abff1b0db6dfc3762f27c3954f230a7933d9ea397a972caac5ed2183ec72716c7, 528'h01c6530fb6b913005f81e156be89b3847701829fbb310d8a4c761212c6d2f8750174f2bf81c238fdde4370fa87de320f57dbed96691af45cb99f3daa865edcdda59e},
  '{235, 1'b1, 512'hb3284200000000930b8b98132341f68419e3262a7f2b8d60cfee7e1e364b36ed4f000bd5fcde187cde7397820b85a174025e4d54d70cbaa80d160fc9cc72d56d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00c009c74ec707252325d78f4e7f14be28f56272be17c0c18c90ad4c07322cef4eea444c8feabf41a213e3e846f8ac8bb7750d49143069cd01877d530bb981f1a85b, 528'h001f1c27ef97f434a8c2ff315dd39d909709775bb3c7588243bdfd8f7c866c49b3369719d5b74a47924bbce57301675e2baadcec438e07e6d532aba664253ab09550},
  '{236, 1'b1, 512'h3bf2ef06000000009638300311c31a5caa29197ef0d079767e66e50824e8d41e5a36f593539a6c0ce102a92493c18061c70eefb94903831d9b8ed3291d1b9829, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01d3b17a34b19d134773988c434a9fb7f22a57dfb4c4bcca031e213e1b9a56db0ecb2f3c54cf9b1b6e5981369652de37337a7a7d7ddb54d67b067bbce01fd7fd2808, 528'h00c90317dfa061122557eb3899939924a8ea3cdd886e0f2e5f2c384b65b1a40de5f00fd9fce889fc313a6a9d5f0a9cd3a7b89b7ba8e97807031f3d1e3f9c103f0a10},
  '{237, 1'b1, 512'hef200f1a5400000000399e032faaf4b3c32d804555abf20471a3a18dc46f3917eb9072220b5d5f994d27b221346631c47eb579d69cc5e438b7e7b963bca9d84f, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00cdca5299e788600a3ca5938d4a4c5f42b5eea3cefc990e67af95a4449aac0ab50e8fc4778efa497223cdca07c0e5a5920110f3a87afaaf265beadbb91c00d13464, 528'h01a92b9a5570b42f91ebc3d8ba272db9241468154783548d3fcfb6ef46c9e037bb6217af0a31ef952c27604629ad5775e7695c63efa138cee8326a51c1b04d0c658f},
  '{238, 1'b1, 512'h7f12580858d000000000055d6877381f726e0a9237d1c012c9840b5b3fbeb6f43027bba37a94ba5fc0dbab436b88d4a7cde6aac151b06214a00cd8fe5f0bdef8, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01660b0ed15d5f63044cb189e1a405bcb591c37217d0e000008614b152665d5bb9353a3826854a8bc6ebed423b15680e4340a00701b17bae24bd399bcff7e0438bfb, 528'h01c47f2f5c6143d2eef063757114aaeb27827b6a8f675d1825dac7f4548cbf78a37eb9621a29e9b14cf61fc6ae49e7e6e15350a4b90a4a897ff69b0c59b69508ebc7},
  '{239, 1'b1, 512'h6b4185d1e7382000000000c86f684e5386df6f2e7e1dab4d1be30ccac1ea33d4e82d455b12857120cfb411b75c8df08758216dcb774dedf1438bd137f831b27d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00364684856c7c02bfb2ad2de603d10883ca93c122d4cebef276467a9b7620fb530e4d05d07c15ab948b9ce7682561307913b64ea6896ece1095dc64369f1a9d5c0d, 528'h009e6db2ff96d9d71150440fd44992656ca118fcaf6bd04499314e8ba61a55a8790aac023ddb68600fbd7ed4cd4decb176e8bd7822ea31d75adcbdaccafcf510c26c},
  '{240, 1'b1, 512'hd40c1a66696b7a6500000000ebb22b0b1f80b394770ad61c5c42ff0584ed4c84a3d185d3c07725f0d3080b451dad86945cc9b0801c01e0b6b8739ff8ec36df22, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01a317e49014f1bf3afc09cc048531010e2144b662cac657e51b32bb432d274a730b535fb2de66fa8ddd26faa3f46e004389d25517c56e7d8a1d39563b0e8c9c215b, 528'h01ad2e1212e1680b660a1c07f54addff575c8c8298e26a14c516f517fb5f966a2b383aa46a483fdbfa72711d60c0f67a2c03d63d2626ffe271e0ce353a4d4b09bd5e},
  '{241, 1'b1, 512'h68481d736990000f3d000000001bc2164f3bf7a43f3c7f23a875b84fcc1d1395c9bc3eec02e9aa7d38f4462d5734ca53f0db4e46498d1b8c9f9f4c92f4fc0532, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01c09b29fc4da04e9b86097bd6d6806aa969ceb37ce52eeac5e9518d27541c3f30c00f113d9dd3b007dae6f381896d43fc6ddfb3fa256a36529b054e416ed6380599, 528'h0113e5622cb1e4c4bb0842f3d396d7e660241116e94e8120a602e3d2952701b1a11415a3d8c503adced160450fd13157ad147d2d65d77449458659350e20a545602e},
  '{242, 1'b1, 512'hcf9bb31b573fa12e7e51000000004b37d8761e5d50f214b30bc2b134bc7e0e30653b8debc737a21392357313d13e08eecfdefd8d37bec92b680a84f5430fb57c, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0078f4a2968460ea8f64a938b3a97c914eb0ccfa94eb08636efee9d5ad8668ce1c9099573abd146df9e7b2ccaaa1a25de903f85962849356a872e88e545babc28974, 528'h00f2729e9593c9fcdf5971b21e367ffdc87aa7520393527c6f68ab512b88b839003c1c9952b04f2dc74010a31071ee20a9fb1c7e1187d04de71b3f4327df128ccd43},
  '{243, 1'b1, 512'ha678a93e12f88e59d6307e00000000bcef462484d98a07578e5106f6b5e6cd1618aa82e3797b4bf519cdc4704616039255cb3f05fc8b93e4a48e2c4cd5333450, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h019faed147a76b65779d0989e1300802844c9ba09f338c5e31a24d9ebf8f0b0b4c21f59d369ac10e315fa2b7605b0f17a9c07cf6ce4c83838e58333a3390142d79d0, 528'h005f4de71fdaced1e8da86efd47ecbdac6a6ffc6d69df71da7ceb5596475cdfecea3d00f074d2de89e0fcc05e3231d531f0d38f2b7c6fe4ecf67a0cdddc21d0867b8},
  '{244, 1'b1, 512'haed2cc5334773206d7170bca0000000081dafcdf0acf2107d7c016b54b1c0ef3663c5ba78277a328ae547ffdf6ef2e385a374d9355022f24dd05ff9b357e5039, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00d0b144350a2128f042bc1a27f6c021dad1ec031be8f1d8304797f9ddcb742974aae209f014980174b9d4e434e3f53247889d2da4b767593179cb4eda47e7996430, 528'h0184d3416dee35ba8807703a91ac927096c10959a05cbffd8103a93a9f20a11537bed7a645f32295e4abce493579caa4e2242060cc4d58b2414870e98b9336795787},
  '{245, 1'b1, 512'hfeac570e6cd1481ff79f34cccc00000000eb127fae412cf598abaa6550b4f5f2e1537dd5c5d6c57b0b52c103ec0340c9e292d0a263d74e44301efe65d505ff9d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0005257a0f45ee2ae5cc30283d23c47c96f6deaa3ac1473e8e8a40eaf61bc4b0ef8bd18d11983f257ec4b1d8d04e76a122b5bbe1d31065159072c58fd9bc3e983768, 528'h0122dba50d0eb71bdbf092a94a7ea280412906e1f849e91dbd5d8158e3fc6cd12e20461b77653e3df2e45b86883f81071b33651ae1b84cc8e7c365ab8d6a36d1cfa6},
  '{246, 1'b1, 512'hbacfc820b1f513e6a157534762b6000000008ba56a4c814c4c12a828e658c8f7d0453900871cece52dca13f4f1df23685d1bd43488e2acdda903b2e0f72b9d64, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h014f624af9d8096fe7a290651d23ab260da64e44b886fef4f3881d0d984d3b387fddcf65b1fa1dbb239028fbab4a1de6ad150cc8a4e4db0a971bb8bcf01c4728ff98, 528'h0105e3b55db0141c06d9854096cc0f73415dd2b85a331da50cfea3bbf648bbf8651f61f2cd09386b62fbb8ce67248683c260894d9ed54d6667ae02978e38ab99320a},
  '{247, 1'b1, 512'hf9f58ffc6e2662f4992e06774f928d0000000084b7ca7f7b6fb750919f466be3366746484849f67645a424ce6009fc560031052d0775f47984d3a4727776b916, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h002c952d7e61e1097cd7f709e62ec486879b380b63791c146b545c064e65b3060250d00af279cf15eade67384b28594db542845fcc6574ef5d8d5bb8a162e0350a00, 528'h0135ac6d1cc05b095fbae28b652fe5386b8689e21a14990236d3ada7ceeb0c12a4f774bff7b81c8d07572b0c7985364c5d31f33271f0ac3a2afb88b46bfeefbaeaa8},
  '{248, 1'b1, 512'h5f6f67fd931001c593ff6f8e5ea8faac00000000ecb4ce9ec81a128cb55bba07a9b186b28f7e787f7bfb7ea32d9047b830a99f2ac4144ee3f6e07ddf00e68646, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h017919eff78225e1937a921f98f5d153cbffa03929819f228ee013f8e59549b04b9867006a8df25a93a6a25dd1d3f540239a8ed14047ea00811da9305ec515ad000d, 528'h011fb873bdae1757801e575c5df62cf82a1881af3cd6ed17dc50edbe6c5fd0f4d31766670b2aa572a9e6547b36142afa8464d0be4bf41930629dc04c85e01b2ee8e2},
  '{249, 1'b1, 512'hdcc948cfcd6f3cd3760d678a643ab0ff010000000095bdd5dd5c0b9579c7c6b0f3e921033117737e31acf8ab117b62ee54a25abdba306c71bb0c3d60097a332c, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h006ac9b370067b13ac2b57f35d6d9b1faa93b9b068ef5ddf8bde3a54024810aa2226560065b0cb7501df96b4756ce1e1fa607f86a942367894a1f7728bd5f22cf177, 528'h008b47a9e1370c9f5bf4677d554c00e9ac3ea7cdfc78836ac53ac710b7f3bff8c2297780c69a9fddb80e03a605e5e48a52e52fd35f41668cd9064886366fda206086},
  '{250, 1'b1, 512'hdfc50d9e551fd99c3ceeeadef83e2fab3f96000000003206a5e2b462805d83d6ef6280540f3bfbb229421d6f5f2794f117259f9dace4f82dd57889a74a0fcce9, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00c4bcfff265cd32442220976ffc7e4ec09181d694696eb89af0cb2d5a2dfc3876deb3c6adea168965200c355c3bff5e47ab17ecc44c8434333280796d3a183449ea, 528'h0062debe91550f8a760eaea309f48483c65a52c7e88a83867c31730cbc6b0a64d4c564bde67e6539af787ecfd18016cde46ddf91740f58f6ea6ec80b173fd1c47ad0},
  '{251, 1'b1, 512'he4edde495afeff435a69e94a6493e4ec2c0b1b000000004c8e512f917698225b0189f732d3deb6d8c1c39b6b59e0701bd7f7605a521891358603454d151d8e7d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0174d744ddc631fcf8202fca0ab10f6d96d3f7552bb2a9ae5ac573634133f61c59a120fedbc39cfb521ab0cd572afbd5147981090d1dcbfe902e03f0c0579967b581, 528'h012f59ca927c4ae331d2f667fcd9ec01b0b5514e2ab5da0561ea614431dc1fcb761c351cd1211092720ebb7074a5128f8019b7c18e048d5ed3573ed61686e9713f72},
  '{252, 1'b1, 512'hdf8f102f7c54ce2cb6ca609ce724818f7621cdc600000000c69bb15b7c33f6b27c75a153b581d47b99de18ccc8105fc3bb697f180112706c5ebfd6fc6c8a6322, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h019a513cfaf871287340d8a51d2f4348ab4096c5fe244b22add38ce433e3178e8ff5b2df0fe74a1ba40fe8341f734c71f9a1177b41035777e2da6b082e0b566690de, 528'h00d0c43eb33a817c3aab30281c593c74517ee84e958b114395ce0b31fcf30bb8f5dfe60dbc7f6f14698977d8e0516a9274a5bd71847057e006fa315fae6922eaaa55},
  '{253, 1'b1, 512'h3e526c3c1f02aa2e007cecd9e02f7dc3d06f361a0c00000000f8e183a89a7218d8183a928d91c6bba47d950bf841396e5fedf9d87f66671deb8d2ebf63e39751, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h013204800efcb40ab09ae4137325a3e8c468edae91880a51616ba61f3ef1f72fd89feb956bfb39818d827468bb4475110a04779fd6bb3def25c61c4ba60889ed0ff7, 528'h00704b7394687698c8841f4875d40e5b3c914f154ccb2b54466ae163ed3410f20d0a07ac5f90c0c31271ec8a524ca2dae4b8bc4f6e1ece173ea907890693c5f2190c},
  '{254, 1'b1, 512'h7a750c1372a8d9b00991182aa031522b94a1a7f4509a00000000baafee68e65ef0a94f7983cfeb9241e0b7d8fd590a0d55b16041eaaabc38e982aaaaf6eb75e6, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0180241cd2e6163158a39599890dabee99c2c86b88accd2b04b5a72874fbdfbde0d18143c4d78e0da1abf3796b238738840d60e34775a8ff810d58a9bb3559a3997c, 528'h00bc396c2ef28b244fb8e004bf5361572ba1fef6fbe081ed1dedba4d9af78deee126599f75a0a9d0f1b1618ded7a0c5e672e40917fdd30582460da3aeb1e9c4477d7},
  '{255, 1'b1, 512'hb8df763eea0cf11e9945dc5667b0147cf8684d618abe1200000000917eeb543a4dddd7217ba71e998bb9c5fd62b57509b7cdb489bc3b64f66a70e4b5c12ffd2e, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01485fc03fcd629fd4c564775ab6969bbc696b5b0f38141b69f86e052e7fe8849a64af2dd37a2adf64672f20bd6f97cd32f0efea51aa22064c5f10a3911177e1979d, 528'h0180fab473ff9d726db6d266541a0bddff8610e4026d26b6c9abf972eaef477d50670bdd3067c9d711a8346e16869147751e89b4ea75bb00ece71300cc3b80cf8899},
  '{256, 1'b1, 512'h88670299bf6b255d331cd40c7154c438fab9fdd2b4319e440000000057a51b1cdea2812fd594a8cdd56b4f5cb069625524bd53a5f304653824d4afbf9bc58d02, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01bea49b150a27026fdf848297b0491019f76abf90f3e6d782e3d3fa6caddb81b7ef58b27f1b2b3f7898889b4e2b6cdda7b5636177a27eb9a67b2055b6f21d262c26, 528'h00dffb13c2d5f746c8573aa444afc8baf8bf881cc4d0fca8169f6cb304f400eb3932666cd3758c437c9cad79abfd89c72a788505763aabdfabf8903ad4a70d9ec9f7},
  '{257, 1'b1, 512'h295422dc27dfac13c79d2028d3daed64c1dcaad525dbbf14a9000000003667b1baf41fd9137fa0bd8c3851590b206aefb6cde62fb4ecc23ae308e540e83a7f09, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01d56bf6f3758f627f470706d1d28c28fbfcad6dc30465cb285a274fc057f791de73ac30baccde044473fa9e3dce6d395eadf98d1f97259bd851a1eb6f3d31d2d756, 528'h0033704b4ad37300a96682569f4f7fea3e14d6e1f65864663f39aa67f40b5c949f198d5de9f2ac2369bbb9111c89b393199537c6c08ed7c02709c733ef7660113d53},
  '{258, 1'b1, 512'h118422376e38638a08705cddcdd319e26fc8a2e6d4a4d1400fb70000000005687b339ec07f51592f6e254c9b7291fa2d0302df9fb2702857e3f69bd4fba01654, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01554035ba84b051d50901c622b98be4de0123a02928dffa7eb13b0403fd5e255f226505e15694956a66a878ff581173d123d1b24eaa85c5fe46d8973a55040ff405, 528'h01b016dd6b5176ad8347eb9802dd7727e06a29db33cc946f809a42f9193040692b0f82ebbd04eff9f099b7f75f8e45e74ac00a51a9cd4f2cbf5f03f4d2bee99c24eb},
  '{259, 1'b1, 512'h5a4801a1f7ef2afbf8e0e76cbd6e07212568cb47638e22e55f8e6c000000003a2aff81ce04258211030942fca855cbc0ef482027b17a7ee523b15483afd91355, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00293e8d6775f3c14183aecc22f608e9013d7b15dad167bb38a1dfef6b373619f1ba2751d77b43f643f68643cfdb5c04a8ed858bfcf3858a681ae93bfc7cd7e31438, 528'h002c7d96db7dbbe347bab9f6f7b88f48cb32ab963248737d2c901b90d64591cbdb0f0ca7a14557f8a50fd80d402f929dad141141f1f0c85d9414b32d1fd4d796e6e7},
  '{260, 1'b1, 512'h057d7524efbce651b92e0a70e4454156e7cd4b696c197c6a064032c100000000768565d4af2019fe3247dba91948292af777f107fdc9c3b47659eaeab26ead77, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00b16a9b3aceece85908125f96f6cb6b1afd0ef04171936b3766f8e43beb340d382084b33439f775a29a83945da8efc4190db1343e87d8c0ffb97aeb3be159d90f59, 528'h00e5c2bbd98e449bd0bb4f75a07f1a88dd63c0602a7660f4acd33937c4913a9c16ba44dc5808892ec88a4255109a7bc5b221c07e6a278888a9712fc2a25b374427e3},
  '{261, 1'b1, 512'h31ccd924b687a2a6b70f4888ea911ea38a686e56e5540ea692ca3174bb00000000246ac69c46506bd8fe924eec33b33ebc9f508d4251c459fdcee3b4c84d4ea3, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h003b47a8ed52f5b0566365313520bc0b6e4e4efb3ea4176ed7a352c4b2f8bffbdb0148ff44f3f13d9e5e31b1cdeae097574aad8bf393c54a5c842e749ee87a74c6b0, 528'h01d3f484e9e224bda9c8f10fbb74bbb62d7a18245707f4eb52f17dde793892c16e4bdf504960fba55da487f542d412b1b833f6f46336118618fcff69469c83963777},
  '{262, 1'b1, 512'hc7b70cc4a55d55342487a4469ad2243ef6d6b69f11604b8c12baa03dd3e10000000014df0db29a9d4d54b26f4047f3e0c739f7a260768b20589254e1235fc590, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0128b8988bfe9287f82ac97be507a544b823e85cc2813b6929e63699cff85a40283076028e7bf8d24330f89adb96bf24a4e183a898e679b36768909574e7d4733d61, 528'h00c18aae44e6801fc2e3d9c7a20ff9d42b46e4a31ca37772f8c46ce65219b195ca23717f816e1fed51e5b6f9a0ca12c3cf81ae7fc9cc6946a88330b2011ddd160930},
  '{263, 1'b1, 512'h1634df8a3271a99f360e3bbdcf789d24bf4bb03e3114ee9f0fa930541f1ae0000000008d976fb74f27eb316ce3a24d92a53833e600c353300f5c4fec6b28c581, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h015edf1fa95b17159f762d68c1736101309e80fe5b2c4415609a5ac0837fe5901f3c2d3d826a43b1f8cd1babf494ffd96cca1267950188a924d4e1bf7f68189f27d3, 528'h002e8697efbbf53adb7cb1b904718fc71eb2561f331c209c50848b5bc50bef77c5c3487d285bfaa3caa14025cbb71bdbaea6911e3610335641d2799c3fd75019f716},
  '{264, 1'b1, 512'h8f90b6a8ecbb870dc24832b1f4719aae2d8eedd7faf97848b08d2b528abf5f44000000008877a6157344e6a9dc43b90c8e2dd7ab9bdc5237c912e094660d0878, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0161f64bbe93fdc0e61134cfd4c453ab740233b436179351aa68a3e38a83400d86ff464d7ceb7a51f541b86eb2f12e32a879b3a29bcb92e08cd50e74f86a0ed52ae9, 528'h008f6fef49ba12ced6696f4f6d24e6c68057a84496d42eede630199e9bd06d91363542a9776bfcd6d77fbae422e80fe466edd2c2c5e1f5cc79bedd1a7becc1a12660},
  '{265, 1'b1, 512'hc0891fc626ef4b106fc00f5c067253f26a2868d09aa2ce029466f353ba525e757100000000a3cee37421995445fae741697659a406394c870d8bdda130080d15, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h013a6faccc1c06cb5dadb2cf083cb94a7181fd5cbf3954fdc430c2691248fcfcd13767e32491f00269b549cae93777ced0f7b069440726adde7605d4038d7b5ea4cc, 528'h007622c9065f4c49a6f8649073dfc6a827b897b6984176b1a09d151b9733a68f6da746c47427cdeb3be075da4a351ab78dd5e472cd98d1586edd6ff2a11c6c169fbb},
  '{266, 1'b1, 512'h76527097fb3945436a30cca60392c170abb7ddf6ddae93e3ff7651d468eb3e14865700000000bd314c31706f8e4d1d853b151f5afe680e13cf2f255b2bb697bb, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01899609e7f7cd2ef14bfbb1cb9ba9283ae11a9346a34bef23b1c249da2e76a7708e0f2f97f819e4e25b0d5227eeb85aa593c3fae9398a7020f61ae1606945d13841, 528'h01b8d5e9c4f030295447106d2b5c80cc2e7d4e36b458a90a08f505df62d2234e59d08187385ba5501049b34e12ec92f7839a18361a52a9a0b6f6a664b118680b53d7},
  '{267, 1'b1, 512'h41d43cb27d4db522756dd682826eee8d0f60163c7f3ce67a39d89d7d89e24818c354ef00000000cab56830cd18f7bb9a7d1b2440fde06ce647518fada2dc988a, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ddc69d1508021eb560db39f3add8a28dd7fbce417e5fa1f4f626705caaad72b634868d01dfc474e926c97927c56ac51f9bdcfd0e7627be35cc300a0cdc083b00d4, 528'h006e862caf9f2df11b0a46104e78865fbbabe30bfac0b1fe7f99badc11746a288c1ff27f6fa2aaba6441bab0372af906eef083ff03ba466b896c9344cd396dd46dbd},
  '{268, 1'b1, 512'hd34ac40ed5ab79a4e5ac1e4081e0e47e4fdedac1555b01ab62a13ac0ae9dbc3c23f799510000000010116f328ad1db0cd68cd1db9e1b34b5a52ebe9b8e372b78, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0117fe2c21f282c7e4a8415e9c53c254514eeeb0adadc771adbc6d21a09add4f17ea0c597469488238be795f2e187fa016d590535b4ff10c62d2246aa17bb013f9ee, 528'h003c9f1590ce7a68fc84c617f478188e71aefe8c74c4b9979b8c9196bcc262205aecce5fd2bb80c360d3e20da20e36c5ab70d810d4ba97d13858199d3a1c9c140c63},
  '{269, 1'b1, 512'h8b5db6db13b1f5e609965dc38215d14ccddf66a9d86505a67cca37f13cc420803c1df80f4700000000b044bda09a83e4331aaff90c4faceea315e467f5fd91d4, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00be6b47254a3cf93e2e276adfb072256404744070d6dec83ef34e3e6c119206422bb275e61fc47053ef7b2af9e33aca8f8b2e4938057070eb6ebbcf82fabb44a5fe, 528'h01061ef80935ff6d0e9f87f3537b639945acf50c5d97d30b4b9c347e3f5f5ec02b15a376ae754d64b2efaa811b3d12a0fff0bc689022025dd2f69f2f4b40dda8687a},
  '{270, 1'b1, 512'hc771e022bc376ffbe1f513bcff11884e790e53878c197014931f6360c517ce8de1c059d091cf000000003c560cc443a6f005ea58917a52ca9bf60163afb16ce8, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0130b6fd7dec5cb6f90a8b54ce7b58c61b013d0aed7c4a26639de80aeac3d9e3388e9f87e1e6419d3f0339af324e1421b5d130317ffd9d8be36500a84bb41d026cea, 528'h0176b460a3eae01d8aa8ccffb0d6cf4d1595aa697c65510a1197b97343c1a6234552ce9d6d318c5f20f48bec0dc311dd62eb40058f3cb22fa958edaf9ddded191a08},
  '{271, 1'b1, 512'hd9cb55a3f1ec161bf6caf0452bd6d6c876b35dd1000eefe18378afaef6280348fd799e624e573a00000000085b3b24635f5c10770090ea935f198728655e236d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00a87de42d827ae1f55d6fab3277c7a9fdfac3af22fe47e52bfee34fa1ee3e765095fff20175becbdc94b4a5ad3a149ea7c1bebf4d45370e6b4404a0437d8fae264f, 528'h01a3c1c5186d8aa491b4623f5765a388930f37bb8f3e1c0db508983585b9090b3aaf22bb846e0fb6d915b5811ac55e4d6cb08f605cb84deb55ab7fba2dde8736b1c4},
  '{272, 1'b1, 512'h0caacc1f43ee27ec7ad5269155a66172ac310d4e202a9b7d3defcfb07ea8da85415ac2b116e665830000000009887d6c7da6cda824528345e14a6675de23988a, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h010e46055d9aa087f1c4b6056319cbf17a0694fe073266a3f30363030e345a4bd461acbd99d1261fc05ef3c9a1c37afba6e21c2d513ea3d4709de5586810d7d29ec6, 528'h00d0c95c7e97a94efb44aa717cd6ebe82de0644e32676d197351f128ee8d2b223ab476d3e66014ecc003081f7040c578b8984628d6ec80733f713e26b2c98cb4ede1},
  '{273, 1'b1, 512'h5d761de2a231df86c0fdd90da20e5811f7bd9bebb3f1966359b8fdf554f79f0bdd32ca06410e70e61100000000ed3d4140a60908e85f7fcbd26dc792bedacbfa, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h012c04d08a7a2d07403aba604ea85ec23a52b52786e7fce04170e867be6146eea75a7180f5d4f3b82a204a3c996811a1e61a3e76ed209c22428b35c51fe60f3bee1e, 528'h016f2feabc25733b0a460463b9933e6e4ae9f4124cd0ad3785c77755dbf0848ec1cfd2ab08b960b556870fa00388d23d9a9fa3112ac3e62a0f342d58fb1f0aa81748},
  '{274, 1'b1, 512'h78adfad2734b7baf32f4e0201bd6c3e9f6c1763cbe35858a0f56466db34dd98a0fbf5b2a71afbcdeebd400000000d3da1a5035406b39aa13c126a3946b6c6a5e, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01ca9532c9daeb80d0dbc07a4138ba62a6bab8c88b9e1e2edf2675132eb97cfb26f4c395f3b9d1d1275694956b34c3ef72cd00bab86777465b9edba29a41b0114c62, 528'h0140eb6dddff253a7ff5b032d82fbd18e481a376fe242f6405b81b57165665c9bfe61e25cd3358245bdfb8de7632de72ed20cdacf384764096c8fe3a376563a348af},
  '{275, 1'b1, 512'hf1d6ef224f72b83a109944afbfb34ae1f70d6e50eee54a91faf8ba0fc062563113d988f2b826c055ecc61e00000000554878a7e761e75fdf1ed2ad2d138b2974, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00d609e1f1cc1adf5889dc6deda441682e760be08932b31592fef3ada143fb4940e4ea75ae519e4fb0769c4fbd33a52b183a21d0bba1ffa3fe50fd11f75c6ac58ff6, 528'h012400cc4ddc24ddcd47a6d639a2abdef29a65d4fe9175f51b316f4bf918bc918879495c572f8e98364e2e1aa0d4d53ad29e803a4470d94dd06a982a1d041bf2b5dd},
  '{276, 1'b1, 512'hb33f308c5b107050cb2e513fabf8b896e52c85852fbe32308bee8b8661121bdac78f52f924cf3d5690ac92d5000000004f0f619e72ec1464166078ba3f508a66, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h003775a7e61bdda9a3a990ba9fde98f9d81d4b03195547bbd0658e1059daa00da9270671b2fada1bbbf13982f87c9f3f26dda5cd4f24de63bceb5fd9390163c58d26, 528'h010a03e4ba08f9e2b6915a6c0b83156b00f59efc5417394c51ca7616b58cf91ab7166d8459eb4eeb0d57146ed6560e173faf354b4390817e0aafb38294df25992cbd},
  '{277, 1'b1, 512'h0392f8c2dc961605c5693d9452731b6a8292ff57d6995aeca0dad3117459668ec7809dc09cf154170fcd624be50000000026e3d92dfdf1a2abd09392468117c9, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h017ab00a30c88faeced3e4a10f9c63785bc29e9af4499466bd8880827cfa580b6171f4a20f36487f7b94592946bca4162faf65872af6bfb1919e6b026c14e51e2740, 528'h01927515f6489e9b7d9cbf61e103295857c8131320217e7a86d3f2fdcb350da5b42c2dbe173fcb025d14da239d7d610de8475914748573429c9590d3594f4fa3aab3},
  '{278, 1'b1, 512'h9dda0539bfe47c75bc00b014dc6046c9db5d7a5723acddaccaf2aac7a9250b732a80cd948409f132d1dd65cfe91600000000d53c76be9f75fc6927f818acdaf7, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h003b2ba1509aea9d42d400400033952a022fe7e00c7ad65c39a2f76d41130aada99c3cdfb9cf44575a2163de29f097beb9bd3aef9334e6fd0813dde2a087f938c5f6, 528'h001afb56087dfd5cb4fff6679a114c340f3a59f6b3e1813373bf3ebe30cb5e8b285a5875d1b5a9120db80f70310201559f89bb1df147961d1ca4fcdb5e8e84cae082},
  '{279, 1'b1, 512'h572e1d736d78c42eed5ffabdfb25b5c7908aa60728ddb3d36a24c285db9ab996433827aca9e23716c3baabbbb4527600000000b9c1a728fdb6f65c10935e9514, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h010efb321a347625343f5126ed8545017d799eb103c75558922eabe44211e8fd834655dc2ec5bee9bb3e44350eb6885e0ab974730222e55f13ad27c066722fecaa25, 528'h00d62e3d7ff9215369aa7da818db302e49033875010b2f9b73d25ca5b9bf2c62ed756686230cd5f4a37c1fa881c97e623919fab827de5995ab456a1fd7ac7b85b1f8},
  '{280, 1'b1, 512'h81b675425e8c528a0a51b23413c8b796411a01b207e0bafc5bd2a46b05237be84abdae1ebd492fca053bf7e3133392720000000086ce63108f1dc5a3b34c575d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h002f778cd552f54da5f567f47e6979872ba130dc0890172bf3b3bb952f03c64bc8783abe9f056d60e1667780f5ea88f59ef33c735d540561a197d31fe34853a60a52, 528'h00bd2816f06372f2e3f2582d53e583e133a551aaec04ddc2fdb7b8131787e73e4295ac28a9604a2402ed5b272cc03be57dd4a7df84d9ee24cb0c2bf124ed927defee},
  '{281, 1'b1, 512'h11c203ef3c8978266a73147233f7c9c9d16108a07847ff587f1e865f28519e7a161664edb56d9e791fba0717124717b3c90000000013c59e26ab63c4a99b871c, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h012a459fffea70d3bfc13e9ea0abb10aae3910df604997cb5e4bb0548abd852abac6b9a32418c3b5ed4e7951ae88eecc0a2f1065caf24c6a814674e95682d9b493f2, 528'h00e2abd05c585e0c213a219a7e7d38b810d252ffea67650d4d1994a41c2ca325bb964920c6c2545381c45ca3e1eca05e00514b366cb0e1e49b8c236d383b260b9cbd},
  '{282, 1'b1, 512'h5de83c97136ff31a90ea5053ff256d522819626ae3734c460ea7681fbd0a94538ed840f3bfbf8055756e761d8149786b8cb000000000f37f36e4d32d46cb9bd1, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h010f2653d94aa28bcbd667a5013f9b283d8487c44d093ee47660329398caa550ca9c9388c7aadeceacac1507e76590afb736adb3583f54f31ae25c9c717ec9f89b5e, 528'h00494448a7ffe4a4eed84b4602781ecef77a23fed116b1b791b8d2e4231b7ca2a7b6f06d132705932d446e61d344714ee24014fa5bb144a96572b3d48d038a55ad68},
  '{283, 1'b1, 512'h4a5e1e8c073ecb2832fe0d0df42a72ce225ea97ce093ed320aaba00cab25ec3e90a6aefaae72ad40273d7309e40582f40a37c1000000000b1e8576da0eda555b, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00c2da48552c39d94f5a45427ae9dcd891b65cca33e624ad2532ffa333666b241d873336fab7bbd7b4c193db4d865cd50f0c1d8cb5c14cf3f089ad42dd43cfff634e, 528'h014f2070dcf860b96a45f2a6061e4ec2a6ad64d7d0e9fbdb25aa93b99941be280f5c70c0e32b6234df545bace7341af94c140c865d44fa8ea7ebe0fe53bda44645df},
  '{284, 1'b1, 512'h9f920bb92b4527d54ff6877b80c81585dc4d3d1e96fce780b030f9f371f8a1b68e2e7a86536acc3ce96737bd5fba0ff669f6b1600000000000b5868a36cfe6c5, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h009bc6e74549b48a1e7c181b179687fb27d6e9acac47ec34b1b8bd044d329320544e4e568e67d17f4cda2f0a3fe303d561a11fc0c981ed9be2fcc6d397a43ad49e10, 528'h00ff295e43fec5b68b00ce8044434bcd17af1ba04a74556353e258d017ba26bed67f458fad5dd8e7d2734d56f59928c2419441a9e8c0573db3586ca056951ca935e0},
  '{285, 1'b1, 512'h99f941e73ab790b224ce0a799133f6b04eb9bcfb2fd0ec84b8e7d5dca6ca50d2b1ae4d31c57e2e54f97f59b6a10d0758cfb3e46500000000909d4fabd9d1962a, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0020963638d0b058494254efce57778ac65e5f23491f7adfa72e4713b7c03946b543c014d9660d855246f308085eeee495cd831b7dbece47aea48e90433bd0fe8184, 528'h0161a4f4977fecae92d4f67e56f3338c7a9b820b5e05db1f28d05d71f7e5f36bc63f6edda4d3c1b2d73bb8a30c4d745b73e634ef574cf47656a372e3eb42cc038850},
  '{286, 1'b1, 512'h202e258cee0bca789ccd4c29f3835362b6f1f53faded0f1d58f4ff768f6202a6de3ee3b922546127fecfdf1c0446605751df9b7fbb000000001a8a11a3e383f3, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01bcc5858597ce8d4dc5ffa6be33f7d804f2f8ef59c5db9301785e0cceb7ed57462f455a465710c7414570c9a35a3100bd15fa40e3ec350d1f75406c2a25885e9d76, 528'h0043757d282fd1d44c253f9a05d8142c29a6d63c0a1f5508431bc9fb9b60a38b7f414e730e0d59b7b709706a67022e1922fe88b182a57443c58bd06a69ee7814bcab},
  '{287, 1'b1, 512'h8c4a184638926ecd8f6ae279181f9171181295757e3eae5b5a0de2fc0281358973a355e4820da4ce0c69db549c72ea007f80ae990565000000009e51983c039c, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01240120b97ea67bcbd0e412d87137a13e347a870a2249375fccf8c004da35e592620774160e7b82aed1f57997fb015a764d014d4be1f389e5499777054576e7bf00, 528'h019f157ec3a2410853274bc4d8e7565e9eaa5dc47d5e515abc86c22fa6dc215482df5c0e2b885f37baef3a6ae83daac930617a5fb37bb03ce40f06fa4ece26cbb11c},
  '{288, 1'b1, 512'h92eabef5ab4296dba863345a2f11c2bc8d32bc02731323a19a88897aa1421f384448516975b6397a8e627fd3cb5a5dd6ee3c50226b18860000000077b18d5c83, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01a7536d55876f8392a6eba18f075118c273015844eb3536c727c004c1bf23067d57e8fe31872f8bf839640e80e06aba3c0a365a268cabc2da96d84550a569f17f9c, 528'h00e840b6a7cba718d91103faa134c2f63763f3b6b91db7ecbd3b10f10171a875712cb9384325411beca9a3aa87aaae3902c282d2dedaa1cbddd40ccf0d29975df22a},
  '{289, 1'b1, 512'h4cb05f07197bd719557dcfbe1edff395550b275100cb073ecb4a0987621f83a5f041996f63fececb77a30cccc5f8067e36f650f7defb611b000000006a949e2d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h013f72be1c331214f45007ff72ce54afce1c910a90e4ff3d176620ff3ca976c2b62d0cdf5d1134290ee97440715531455dc29818828094d366f959e1adc7d7e98ea4, 528'h01e80ac38ba69f3e53116e5432fbdb3b1e7ea1b43e5f86d1c0e3d1c469442dbb406ffe524f0685f71e811d94a9efa9ed38ccd9213f983983035f2add0b8f2fa4ae23},
  '{290, 1'b1, 512'he744eaf4e9c4c17549ca3907721df98de95b69d07d56eef509d4740a3cb142bc61b6c4d108676526d5a77188977d924dc9a8adf6c01adc35d6000000007f3077, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01aceaa6d567ddb39ba52d297e60e4a814c9b476cab568c09d8ace878d846218dd2b5d2a2461f0d5a56c12f0bd803e3253dc5b387b94e86589cb1d0cb809c7071125, 528'h01b1fb021b10b593cf9e793cf22a88bde9a4b92f9e218094f270b093e8c6c95aced43d097bfa3354e6b98d195c599c2e6f13351c63c28967e08b7e497e120665c663},
  '{291, 1'b1, 512'h4fbf285c9be6083627ef151df0d2c5fb00b6edcfc44216a30467a4fe268214ab66dd9be898bea57b48f6499d09d4beddb7c9e8bd813fe7c1cacb0000000054f2, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00f6ffb5dd786326041e74564b719d38924a28329868177c13463cff90c4b09d3d2dbc011281cc78aa0e5e8656123bc50605601a547bb4b1761f852a120ea46df9df, 528'h01a407fdd445614a16a5ebd4ba075c6c1d7564f3cfd477d6b2620abf18a5bf78311282ea45b9bff813f24c3c7854e6091c8055144f9592fbf2e456421a41c555d7a9},
  '{292, 1'b1, 512'he698cebca57a541614e179f28ba51cf82fa0fb4300f81df5fe22b635eb4441b496a36ad280999f503edded3ae1cab1700758b5ae80ce33dbf25c7300000000e9, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01a15af4d5ca3deadecd75ec1baec31c8d43fbc889466475e6c23106db4e63ab69003f56d819ddfc5a673c8289f9e6df806b07af57a2541af694e6489734c8eec837, 528'h0069c35433a3217fcd738a65b7da9e81cd81f04f0ef060050b9c843e9e808d8b8175f3adaefa105d215ea9a46bf415fe2ac180958fcdd878d54f8d19d23e11b76d1a},
  '{293, 1'b1, 512'h43f5ecee4c9b5bcf2497d9753beb1eca8a01c143f8b50518e83bc7f3f62d049b03430a6dbc9236d54b7ef5475a232e3de9160e9649e3c8f46d2f1f7900000000, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00ba899f94841db6c33b850867c8906b436be3853640dbfc863197fa1e5a55ce25240f2be498b9bdcfc0a89dbdca192d8f84ca3c44e5e0ee6f83e7900e085e1bd481, 528'h0086e6d558de8d8f014a85cb4a5f6908627e7a1acd70581d9d9c7d14df44d437aa09e5a10a0b760e98d46731f2512ca1b0240c602b5f0a2030485e34de9c6cd08e7e},
  '{294, 1'b1, 512'hffffffff4fbe152fff953f198736b155220dfe633b6fc7aa5bb392cb96cde9fc658b17828d0d04ece0f6e35ed6bbf357b86665cac7735a3b9c85c038d4a85019, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h008eb5c92dbf5e00888b85e6bf6617017e97c04ae950dd731856b9dfb20e0c0e5c54284f411231fed1d071b321f78618d2a75c139663fb9db3435214cbac5a0dcb4f, 528'h01da0dd29d4728fe6331c8e2ade5045b1237664aed157db2a6cbdeaf5abea81324e28920a1c49c334b1226441f88e1a7f2c7e01d63e950d4378f08973db16b2e6161},
  '{295, 1'b1, 512'h47ffffffffa19c2322e79638701c393ec0df74b5d27fb9ea7cc3e3dc8badffcac83dd8c409a22c2d7a64b5693f153f60264487aabe5df546115cf2eaae415ac0, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0130779f943df098ddb5315cdca4b731c83472d589f4ba4d32c172faf6b3a9e4154c0517fcc5c432eb269b0152297f6df490ece59496bea8047e2f32d0b5f91e85ef, 528'h00c9eb0b56273114ce2e553341247da86b813bfd65f143a5562bb1c874ff970523836bcdf390dc196e67dd75cd28112ef74afd51b1fb35333be0505a012efebd4e22},
  '{296, 1'b1, 512'h391dffffffff5a981c0576acae266e7b35ecdfeddfeb6db903e9f4eab200dba039b146517f0c5b418d096addeab6d0962a6f77c2a2a552748b788c07796553e5, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00593f0132f7b5c282355978a2cba73fd3bd5ce3272066d4ad9bd8bd8b3e2be0990071b3509ea445dd155cf97e294e2b8d1355809d880e10700eeab0eb8ebbaa4f09, 528'h0107eb3d5ed75cbb9bcb9278f2266c14c57cf703cbd8f7c7de45c51f0f3baf1dff6bb92f1cbf89ba649677bcdca776fc57f587ce714e2e43e6cc523f0d0a286d38fb},
  '{297, 1'b1, 512'h8c8ed3ffffffffd5bc0cf4859c831b89860c28ba17ff5a259b6982325be66498c4ac3119da331db0976678878c73473aec528a7107d0d9b1a17dacb9a9237b1f, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h016ded17fad10f945e3d953b4fd3b72898c370f15164bb7712673385c10bf3929bea293e08bfc30029a465138ad47abe604df807b31707fef55adf3e104920038e3b, 528'h00b76b212d74e4b6eb994d926e9e796975235fad90e339a21a329e6eed3fe96b6d3c0d5426e8464c4a9ed5cbe08eeb5e490f72e9e0406c0d76ad076b476d07c0144a},
  '{298, 1'b1, 512'h531341a3ffffffff263c81971e877fd7cd8308b0d536d7fa3c88e3beaad332ef664f76387e4c43dee6c0a06423b18d1b1772f65acb4f9b672b97a648cdd25929, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01f8624ffa5a6aa8d9d04ed1c2272ea55f5271ca2cfc9aa6a3778a0b8a230f611e5d65af18d8251a0cc4ace663878c33205239ee7e8388cc0a040ea51515072e3f61, 528'h002c1e61197229f40e840ea37325f3bd87a6cd32d080bd61bbde4b072cf7a0c8a89d402cd9235c26f19a084ddceb1cc0bae4006251ccbe10de3954e85a8c5efaf6cc},
  '{299, 1'b1, 512'h2639a8ec01ffffffffb54d98af88ba2ae383d69bee2f5fadda599d58796fc766130e3fb8f4ec1afceb8a1c1faa3ad305a0fdd65796adf8ac579c1306d5f0195d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h012b01c6601ceca9e58e8abb85d1f6663df70cee761a756b77e45294f09ae609a6b76cfcd67f60e47a3494cb85511e33d92a8d297a1b89e9a9038c0c5b78c3a3d4ca, 528'h010ef5d2fab59bd42e2e92a2fca7a975b959dfb372519330defc8fa8954bfcfb397ba939edb6a944a2ce9f6fafbfcda6092cddf628801f6dd8cd40cad4d809d5c1bf},
  '{300, 1'b1, 512'hd9753a5a8b1dffffffffcac9aa24c9d687a2088ed837789e72d457d0bc67f54860087c3f0509744e0b461f88893e2de6c757705670006c9e9e8c4c3757fcb160, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01c54a330b9dc47eb88dbf60c9ee49f2c7518c0a78baf642c74105fe283fa4c357ff22931ef42f92d16d6a0b806ef718539d21cad71955a530e21cab49a56f561673, 528'h01c2cc32c5a4d335c48d0cbb0407fb7e4729c57251afbf9534c5309b94e6aae13614a1f2514252f48cc7f143ee761782f8dcebf2fb490e08fdeaf570a7ed9d287da2},
  '{301, 1'b1, 512'h9a6bf9edc61a22ffffffff703f4706318ef947658ec44c90cc1630c916924f1635efd88bcb900db41dad160ea33f8176397bb8593e19199207ca7d57bbd28305, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01467b4511b9d6601da3557b8ed432c14a80e5999847be136c756a88dd5134689b5ab70d0a2e8fd8d6141e2b143282f98afb93b7e17609522dd9e64c9e4a31c7c34f, 528'h00f50ee66a1dfbf86167ba5968d4ee3506a7cffe0f521c1bf830d0867241e345d319e77eeca45858bb3062acbf8d100bc6bfd3127d57a7e91a8199e05052b8ccf304},
  '{302, 1'b1, 512'h4c18a4947b15af08ffffffffb9de1de3873b4c26280b1286a51715dcfd1242208ad49b2aad0864d5a4529e4a653d7a6355b7c1747fa9d876159d43806661395e, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h007af90f6227750f917d65b1c60200c755158bb783a479be6877c59ed89ff595fea3f3a4137591aab23826ed385bd6156277364b5d603ca272259083e6e9ab5db3f9, 528'h0070842eb62c894935b82da15ca611d9d754ef57859e0c912c0358d0820f4940cdf5360f116a7547a81bf65617f182e597eb1007e26c62838487ca021c3829a590db},
  '{303, 1'b1, 512'h6e50953fea8dfead2fffffffff824e02147d010595358c98ec376055cb9ddc1dfe6d3874cf38e8a98ef0664fd3b10605bc14506eb7e46460c9db81b10e2f6730, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00b0169e68062caa79f99ec0c72d83c4d0fc2a1c818665cfed1aba3e684392b9a95afb82ddd1de49e3fc3cb3889b4f5a86a7bdf944361db2cfa57021a7643fcfce95, 528'h0115ec784e042436892c6cc1bede0f4b7b6eb24b300b1f0c674999a6da816dbefb2d53f90b0dedb962a085e5209fcea50311130800d2a9249d279c7bde2f88622512},
  '{304, 1'b1, 512'h1539fd34220ed16ae0b8ffffffff88a04bebde47a3a94f1b86bc687c2ce7648caa7d42ac8693b5704e401b7c9f4864bbafe3bcf761d862739eaee02516a0d707, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01de4ed1ee81d5cffcf8256a06858cba5eb925ee68e3ed848ac98071b6e30c3b44b102a2de8117cce5b4f9e42603225e0dbcb3fcc171d1492e7ed8bcb6ec286c7de0, 528'h00fd1e93bbc8b8adeb7864a2bf8e29d6f9c0966fe3d543525bf268b57cd6fa8852bfe0d2750726d5445560f2fc211aa7859dd3ee10078ef907e49cd64326b397e01c},
  '{305, 1'b1, 512'h69e3c78c7125bdee7184d6ffffffff274929ae7dcfc4692b84880a518de1790a758005ef7d4e29377cd891eb08e9fda55ac99a11b4dc9a15ceaf8887ae941fd7, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fcafa62ee6275443d7277fc46e4c30b4db845ba45b5d6b54faf47bbf921f825f6fd0f23a38c0c7f4debc33add282afad1154c8707b6e18cd65adcb07d32915b462, 528'h0087a27b2bf3c35d18fd397e0cd7159516cf563b98441e030bfde93ceacd2c4e41228b7b33443ef0a351ce553d6d1d71c12092df796276175cd779b8090c4958b391},
  '{306, 1'b1, 512'hc3b630a45b21b937bf78ef4affffffffad33da42317364a1090ed4446da7738caefc807ed99c92f85a6f6ba946f99284d4b9793896bc5e0b6f93cf1b09b35a6d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0078989628acfba86d4bf28beeb9f44001fb8f2d8e245320a19efdede31eae3ec8b496faec30c85e8f63f8ae06046fe1d1575321fa04953e460f6b1386dd5df94edb, 528'h012aba3349732e21a5bb27d7d6facd8c7688b9d0d0271d6a077f9d6d82db45b5456b767f4b9f1a80f487031f9c0b3ea833c63fdf9c6a25e6b424c19c2e55305d7a0f},
  '{307, 1'b1, 512'h14f3b0fc1795c9d400d904ea0affffffffeabaaa40c2f532e33f6c61620d23188712a838f9bd1502b2a5c321117ed6007ccb48b375c581fadf340b0d7edcac93, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0014a5a46a3ba415f6e8c566ca1b15fa2055649687b1a9fc84cc0fa8631296898fe014e0d45927e4271396baa4cfb3675669b16e76c339db3c0edaf61337e8bebe91, 528'h01fb313129757f76754b60fdb1e4077f9fe3dd62c8bce52190cfeb9c03021cc92f6d7d1302b8a84733486bf769ae94d3db4b60b6df28fed481d3d7c510299f0c319f},
  '{308, 1'b1, 512'h386b3f08bc91c7e18354f3d46de4ffffffffbf492f2bf174abad52337a99f29dda6891d96f85efb667480bcad7d2482ef7f32a314b4dd39576ef560bf01fefa0, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h008a3250eb5f28b598c4a42890d25f6af84082d4376f84f1717e5112a76623e6fe0d207c39463d20bb86341bc26c9f68bcdf794671a01f90465025f87a8c52137edf, 528'h001ddd317f6622d9b032223f76765ba6c9116ae4b43a1bd357bc9db6fa62f0867dc5d8f781f08c1cbd49b4424fe8c22cfd1dcd07cfde7b3598342442589825aa67f7},
  '{309, 1'b1, 512'hcd86d593a60faa34608d5bcdb2e878fffffffff06003c116f812eecd35fc6f3cccc1dee24c5cb89cfe9d41b0defa4e5d16b1d9aa4897e6efc838a8a6dd5f22aa, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0060ee161741d5cb2dd0ff2cf9924aca0376b1544681627a31688e4d8b3b63a01adbb417ee113b9ba8d4d13b7b4e1b14b51a24dbc3f099b068d916aa94862ee081b4, 528'h015caff8d30141e1c163e3ec62b7e14874da624a6d8e0252d8e829860e5a49d3732321b625262e5c9b1ef348c3e7cbb1de8227513f320637866785e97e1931d35ccb},
  '{310, 1'b1, 512'h7939a3e06bee091634b535adc98afd56ffffffffeb0206c5b2cf892d2c8fbb5a2e105567cdc4447b476525488611a085b870e498a13b891cfb9a66ad725273af, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00a1ef8229db9f45da38ae3b6d601110611e209878bbd03ac2a6de65e8402957c669a115e3f02d085fe2d031c61324b77052ab346b4b1a437b58062fb36f9d56cf45, 528'h00cc5c0a3b68970279ae16880f6ca579d0171a827e99a46aa82b9242dcc09cb0b22a44ebcfca84293e6d21aeea492f00ba3157c5b6e2e4caea6a1c09c824720552f2},
  '{311, 1'b1, 512'h180c134c29d50916f2c3b32bf43382eeb0ffffffff6178b5edf0856813b75ccbb537c57758d3e55c190bd8e648a79c5bc6a62e45f2f037aeace1733bb7260707, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h005aa0c8a378c4e02bcc2f56c2c365ccee424e2973c28f0daae8f4c3f0d90b421fefd456e749087e0c667c2a7147bc67b90c696244f216b4d9d7418eadc7d06ef1d2, 528'h01e28914bd341f526b041128f2d251131d8b2c65847e541d65adca3442962cddb2a71c64fae39fdd56e41686ad632f99c6038d8de0b3aac4045e0a961efdbf4c6a22},
  '{312, 1'b1, 512'hf2694ba9c9a0d83faff7ff2f06f0495682e8ffffffff1d5cf19e626efbbb1425dd286e93044edf262236a46a82638145b4d15c18aa6e1edc919e22bff3a9c5aa, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h005a05f5366c8b8be28654bc39a6671d1b1593495e445c07c995c3be3e168ffdec92e44288802fd455007f8746570d93b5683e4d40e9d9e59de539f0e62bc40d92bc, 528'h0187a47d8f70adcc5e10267b8fec89d7011d9985427645aed19a8efa2d1189b469cb7aab1998e0c1d2fcac5a5054d79d2ec1c9a00b183dc9af20f555a1140be2dcef},
  '{313, 1'b1, 512'haa2db4394e6e52a9f0485ea08186ed648a109affffffff19fae34ae6524a6abf956c07617b15896bd3dff11cdaed4f9a2769cb4dad0b0e007b66c06fda3f256b, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01e213bcb8b960b1296ae176993b2449bae556b6d90df2f07fb08ad8fd60e3b7fe6c73f9c8a7364417611d60119c550261c54bbca8d61e264130ab90187e27d22dbd, 528'h0034f519382cfacfd07b0a6f3aca117c13d2be725d2f9ee4e5f88739c99121e63ed7358046bfb1575fc73e1ede8339e46c5139843e52e9184bb8c579061a154a0b8f},
  '{314, 1'b1, 512'h59ce78a87d80e90e1e6b70def3179e12e78cd5f0ffffffff11eee1f43a7030f096c301beb60d1fc2be04d27aaec7c385fb9aadcd6fa37cbea40783569080dffd, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00ed11ac7efb1f29ee64108a5e2606fa9af3bbc12d1a952e47240d5236df64f5b2b77a0f7a0a73d30d0708b5b23ac6d584bf6997d8851623793655dee8774549b829, 528'h01e1602a2cae7d3212df47eebd12e2fe404851201101bbde702be9d74d040ed998e79a09ebf6d055f94473b1f8d87c99aa165bdaf0a5f270d46caabb8e88bfa54103},
  '{315, 1'b1, 512'h5d07345f237708f45b49a7286977f331a27c8cc58bffffffff492a29a714f16596215046376e8d35cebaaa06b73f14ec0731a0607ab89c4edee5ad7f575c93af, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0007123c45e6e9338bc9fe225cdd96c5ab36cad5c06163f44f6bd903c7594e8068ba9bc89f652ec31b6e1298766b246c1f10877f1e3ec9829b0937b8d36e3c1ab2b5, 528'h01688bbaeb188b5047be6e8023b14fb121eb1451dcb19f814f5f4dca55ff95128011e3bae505a4d22166d00cb7cf14130590335ee923dc5db3e736832a128a067aa4},
  '{316, 1'b1, 512'ha6d55690f7fe8dc6a67ac00e5f136dab1f6855b53643ffffffff2585eedbf8e7c3db326f7fed8c48851376d7b1a34dfd79aa6837d19b05becbe8b8d122d1baf7, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01264e3cc4fb802aa221d0787cd0cdf44eb6568982a00a6639f15238af36e894b14f45f06f8c2180fdeaaac77f674e056d1928cbbdfc4b2ceca0b35345ca07bfff7f, 528'h005c2dedee6b3aa096fc47ba0991a077ef4d5df20d8eff1bf8354412b171f08a98cea1704c8189a7951b0e7a8270ccb285b8db8e35285ed926b19c1eef07fdc05ee5},
  '{317, 1'b1, 512'hd42f5eb7f42a9dd25a5d9513de8b6ccd5bbbd029263799ffffffff3baff5bcc111d8fb4f14fc4aac37a1dc5633df840644aeb69aa87f390c090e6730bade402c, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00ca3814747888751794b0488955e2aee07e5fab4b9872074aa7432698e7c83b8079773734df1bc752548a218fa59a362e0657b77ae7798ef4a7a3873256ea59ec67, 528'h015df8f1f16611c960d56647424b97936c8a06f62dc3a95d66bf4aa378d7a9e17d2afb53565780025927e6928f5313428f1d6708339787c8f460ba18457d4c0f521f},
  '{318, 1'b1, 512'hbf0fafaf135ee4e03b991ef87e6e9377150ae255e043de57ffffffff10002deb92f4bf4c1770933d3137b0165ebcf81c8c3387c21457e0fe0c39c7c7947837b9, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h017ba871aee34a893c4ded7a2a546da0d6867d428497b80fca7eea6e51b73d6411aff7609743e6242b6d4d3736ddcc9ee1aa12c8b62de5382e5c33d1fc4853e3e47d, 528'h005feb9d9f8fdd44622e4f9effe73fd9b467d355fd6b8de205527f722ee2f5a15eebd59ccdd7b57da26cf953f78886db5a6e5bdd0d56c9bd47ba2271f77687a64b63},
  '{319, 1'b1, 512'he0dff3b5ebca4c971f1da5a6726d24519e4ca71f45a548d85fffffffff415d9ea4bcfbe4749c275d6594e8ca8b76166fc90eaf2d9f466b0f0a5ed8c14eef030b, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01840793684765410baf26b66cbcf7c36658d6c18a2f750c1225520e9f3a7c1b890583f321d4e48752c3b3116dfef733ee386c52a53402acea77cfad1db9380110e6, 528'h01b51985a306fcdbe3692181106d7d6308873912d003946992098bc98b4261fd78869ed8218849459780b6079f6899a47fcb9ea4874d1c08fab82c6f1e9c9aaae245},
  '{320, 1'b1, 512'hd9a9dae1785ef8a49d7c81b0637471693412a29484ea1cc780d5ffffffffb70ab50279ba56f6576dd87ea0cc08ed51afd395238936b4aef7284700c8d5aa9f05, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h012276720b2725ba556d06be39cd16ca0a0351d8f530913c4f0cfb71fdda74b83f02febddc8da0a1f0f910d37d3f5332c027d7bd4c38fd08ebc770bf125207864954, 528'h00637e70b06045a86e2f329f907e079a785d7f8649541860322fb8b64b9736363f90156b9a5532d808cf2af33b87ff970c02e648dc4f1c90ff0704028ec2c2d9a82d},
  '{321, 1'b1, 512'h75c7b98cfddf04426dda027ad897cd5ba9d5318c27288ec0f6fb67ffffffffb744ccbcda470681f3689c70425ce514d035e05dd133da5c2a104980f4ffb91014, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h007aade608b22c77245734fc5c4be8737ba24dc2ed4321b58124ae46a77ea7befaa5bcf166cb966aad007911623af10925a324bc3c6d06f24d0e2e7b2c7b8468b8ee, 528'h01e9913a412300b3980719148de0bb03826184aabd58f19659aa8ca18045f36c73c97df3d12b921de510ffa96ceac5454b801c86c55a06b2d771fa77bca784332c39},
  '{322, 1'b1, 512'hccfcfe85e6d12e377ff1bec515ce149719d86cf3591b3dd8d4344022ffffffff60380790c2be6a944f31e63ee7b421a42ec5ab43f84f05aadc5ae5c42a6455b9, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01eefc7b6c1468ffa7d60b8408bd44c64a3ffaff298168c5016c6f504031867ea14ae48c661b8124418b4ed6ccc32df6bac6d0a485b1990236e15676268b7868d276, 528'h00515d48436afffdb65caed737116a861974b734bd1903e37dbbc231a9db37464ed762e364cac8b32f1546d6de37979fa05f8b80159a0f747d9470291af6569d6d94},
  '{323, 1'b1, 512'hc445da85686a33c8af5997da14f197df87bc3ff9f277b46831c87f8147ffffffff0970446a79a2c801e1a6f9c03509ae9b782a31b3b15dec03f5789a8345e14a, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01271b912ca055040c227955df729757654aa9bbdb73c61ba14155220e4e7132319f6fb0ee94f2fbe160738f1dce2ad690845c38d962db4fda1598e93270da84a2bb, 528'h00b8907f041c3b19b9234ab555d0b48325b0cd330889a53276a1e913bab892b9c05cfa889005b14ee2730220746aecf12af911c5baea4be377ee76c0eeaf47b7a712},
  '{324, 1'b1, 512'h6a94c0cd0809f1ee1c23039f735f24a0a006a0504c295289507a9dc93e34ffffffffd7127f6a21cd1ec975e05b1a8d78144da6293f4440723e7d6062dae06a1b, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h016a813db0f75f9047fb11f3e19fc1688c29328a54f56ae30c1c9d9378537bfc40c5719d084e49a3b4aea255f5b7f6cc775492b5371e6b67b2d6abd5743e10fac709, 528'h01c258ffd830151bfd41ccdabb86b24af846612788b361c196d24e997ccf3f17d4452f63d32851a483072e6908095e5c49bbc241a0417749b097bc1ca0e4d127779b},
  '{325, 1'b1, 512'h31599cefc10a3c6d549bab5b19bb49d01fad30283d27c8a4905d18cf61e045fffffffff3efa7e2362af0fc827c4bf245dcd58374b350097d26ac996598012290, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00156a04c22ea5bdb7871124f1117301d781113ac4c9d4da05fea536e983d9261d25dc97006f8c78de23c788718557cf6f98863994af2086f0be3e8aa8812dc3a11d, 528'h00ffca96b04c56a4a6ce5d22b36e44d3b974d520e7f7c0f9d69034f9e59e0bbdc43236b3e4bfb0f6bde8802cc5cd6022cff166f4c488d64f38d44e3c563da31cf6fe},
  '{326, 1'b1, 512'hefe7f8f35a94b65eb3a9299658db8b8256f29f2df969035fe5769c11e85c9b7bffffffff61e57fc3e05c9a1eaf760ce1b13dc6ddc5516048677e1fcd420a6427, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h010913540ad73ceef7314d1758264e1d1525a371a7b9b3086971599a6b749be4d6ba69269b089508f6500dd925aa89a7c7cb7185e0cca7d2ee5664f22845d961e317, 528'h0135256c79ea5e5768fb3a55e2899b12219b8f68953ccd98c710b6a13de0f59786f4331845e65c7dd6340023a5e280206ca31416058f395fff4bb5de411ff66fc018},
  '{327, 1'b1, 512'hc5c3daa9bce3e7422af1de2fdc992b34f5c8ef3fd448b45f2426e1677feaa86aa3ffffffff6e9d87ba471035c9beb5d2c94f3bb0dfb4c48298a8615840c621a6, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01b5051ca0dd3b20df7d8c5b92cb42b8a204f92fb4e58c612f43d3800de8c0683c427e832ce622156747052b81bfbf6ed5fa177b6d47858ec8478f6c9ca7948fd511, 528'h01fe5710fac0e9d3e2b3b83081b28b194b822d0c13397bf1516140cbe3faa52e908848f69789a741b9cd54d703a94577fa813e2f2c75834807401ca010fde5328317},
  '{328, 1'b1, 512'he36dcaffe4916e59e41b560c2961fba82290150d1b262323c674311ef6c87564c8aaffffffff573ce47a2b2f25bd4f6468ef2788ede75cd3b7293ad2bdb46617, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h008d3c8f8e7ab74d49e16a4c7db3a393fa9567777e373313667f9ce32b1b5e648debffedfd2ff5345ca1b8154c18c8b883957d911e41336285f86261c3ee225fdedd, 528'h003c51b84c2c9a3feb76a6518634b6f09c0dde8a9d08dec0b3d66135cc1bdb0a80fd69636104af69de8f4062646b29fa3af685ec82704cef706a18c59ca7eca0fb56},
  '{329, 1'b1, 512'h3f4f00f697d80c258cbcaaeea0f4fa499e0675441a078d32627378ae08c27dc9e8b60bffffffff59976ce86a303743b716e53422d7a17166a185fac1b7722d2f, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01195625a64ac11c4fc1fc479ef80430eb85c1af77f8a197a17e009569ef6c41ac6f35850755379f478d8928b154e3baaa29e92b481ac04dc72f3728b4f088ff37dc, 528'h000d55c7067877dd1302fdc6bb69b7b7c024e4cf3a0e924102d744ac52366d9d76d5855d3da228c4b67bc7bc4b2a14e7999962cc9bbdc517fc24a823abf584b8f56e},
  '{330, 1'b1, 512'h21b10973b98ea1dfd2b0d7bfe4adf9d4e8616759177daeef38d7aef0d95d226ec8e1da39ffffffff43f8e40342757a93e72541afd7a58ea2205891c13c72a8e4, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0026eb68bc0fb7664c35bf5762cd532dce33b0e396e97d6f4143dc6e1e766c836e27c069da9ea1e74e0b03d030cf8a81490508c1c728f86e59282df94de8d8a0dcaf, 528'h00a9fb584b712986f19ab7568693df278cafa43272dba400ff333cf48b5556e6e78353a665605c70b6fd0f18f30b850e1a47cda42c4c924bca80102e6793be9a8698},
  '{331, 1'b1, 512'h3be3c1c0f8b8f6b9c476455ceee9edbf99283f1eab4a28ace9494eae8da166e4aa1d5def8affffffff3d69a06db8c19c0984bdd10df6ede19e4214183d3b0762, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00f3d34e36f9754dfa8eafab160ca96d91c7f4f388ec82ac33784026bb6c6a035719eaeec3ee511fffb22dd5d6ab819e6c6387192d6c3a6e9249ead565157e323f62, 528'h01b5786b1d662d26fe9f69c370d2bc18882abef693c8f17100a02725de7c9f03602fd53a9208b573b3b7b0b66db971767bde835f9e8f42ada201e7b7391b86fe0294},
  '{332, 1'b1, 512'h14a2049293367e5ace79214bfae58e1007b4977ba9dbd787dd703160651e580fc6de8759ef1affffffff483224ed924c7a2906cccf6b3b39e1af044f2a7047fa, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00e69c833b604075e9b28a2ff73a56a32e1a247ef9ae01e7a0e471f6015c2b86eb864c281c8c93d2acf5653ad05bafab2f58027f37513eb8569f50bd475e770e9a81, 528'h00b9c9d6ce09b53025bfcaa7d172ae41a9b636aa4b80a930931fc99e5e2aa23306f19dc57399b0431e72440a1f4ec7d5ca902f0f7b81c91de85e469f992fdfd4c52e},
  '{333, 1'b1, 512'h745beae01e0b877f882a42a6339b12080d956dfd5fa03fc87f6c99096ae69833fab59c416b092afffffffff5deea8d387d1ecabbcedd6c2334cf7eaa7aa55d84, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01c6b8b5cf3c4dd3d62391f18e97eef3aa6ace0ae2c6fc97a561cb8e49c087dbcf8135fa433b566b3385cb57202f1b12164fe62765ef73b72a94e7a57870989a4981, 528'h0185944434b83a0d0fb4bcdce8ddaadb30a1e440815e7674562df9c8bf711222208cc346b9665d90abedb437912391505dd5d26f0178e7c063790f5518f47d1b05c7},
  '{334, 1'b1, 512'hc09dc1025bb9bfa3ef093eb420b7712374f3164db871d4cb44b8ebbeec2d5b415a73427419c5e399ffffffffb45643293f60ae63fb9ff87c56cb45252c8c7c29, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h009f351a41d5375b8993e90b8d8a65bf01d52d14aba1dbe49cbb4ea823804f2b533e0c167903c8bbc593297c18f309798a544787d598074cbf56ef0e5022520912ad, 528'h01b892740a57204186bd5f434f72d1534b4289f8f7114cb7b1c9cf4541d754f314448cc32deaf35608263488fdc7596f7481ec098b36f8e440829194becc746c77f5},
  '{335, 1'b1, 512'h5f9b29b201a8f63acd7387dd71844b5ee67ca50c5a76a2b273a80d167abbdb6727992779f49b848976fffffffff2d0eab3e1c8f8be0d76338c7e8c92174b32c9, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01fe24ea831199e31cc68ef23980c4babd3773040870af8823a19708bd0229adc1ce99d02e4d95224101e3e974236f54df86051fa1e9fd21380432633b2495ab782a, 528'h000efd1f2a281f967e7b09d721581356a714c499f9b14f781992eb9ae7a19f6825045fdc6d9d763f44e1e7c91480a678a1d8ecf6d66e76cea3505f65ff78cff15cbd},
  '{336, 1'b1, 512'ha76f6918ab70eb9171fdaecc8add5917f130dafbb7077543007be1aa2cd3e446114f1fed5989c6275e0fffffffffd7f5a47bd23e9cd47f4572a1d1146b38972f, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h014c6ee9de0a2a0b60c981831e0acd6636b46ae134fedce61b0488112663b24e1d7e74e227fea883d26b68f21e4135ba0e2069bbe0d9c6433c3908fd5b00182894b0, 528'h006a180a493182c6bc2a09d7e17ff5d62015293f1e8ae205a16fa09042b0a9af6794cb377f4b8b1175fcee5137c234900f735c484feb7da4cbb405cf9e5370fe4f49},
  '{337, 1'b1, 512'h1694c34168745c74ab9fe8224e6058e045c73458f7e43e3884e3ed466f716a7406be99e0ef57710a1cac21ffffffffd497d0337e572f1afbc8b6b4f41a873e22, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01044a45853ada17ca761acc7df6d1d380252cb0fa66124d9278a5ed8a4a60453bc71de1dbe32b0261165948823c461c7c1eb1714ec1dbf66fd602c7a47446d1dae1, 528'h00f8b27f7c71e37e4b440d2c86f1c1d50bf7c53d3878ed27e7bcfbeb902f769f86d6c3e8820b99f890050f0dbebd2132e84626c5b16a8c7ffffc3a30ace69dd15a11},
  '{338, 1'b1, 512'h3c28cf3e9527af87b483e6261fe32cee8e67cbc04b983566b27f8419a932186bce21c021eb58c8ecb0b707d9ffffffff035e36909fbfd832447041be74d2ab4d, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00676a381b18d05207cddd73b44e4dd71449985c0fa7de1fff43ca5155139a1a09e5e3fd754d86ebbe32f6609f6e906d48d24790e494343c61faa90bfdaa4f49fdc7, 528'h00fbc1c891bf6e368fccad51cc9b2c29e8e92b658e88c0d23285af269aff6702a55a0ab16807e5523b6637bbb004727f6f55c51ad4cec8c924f9c1feb24601aeddef},
  '{339, 1'b1, 512'hea6682cf1dadc5f218d6530a15452aaee8857a4318ef3da3cab58358a2e5d0f8fde22dc704453fb8056d224426ffffffff4335e1ab7e6e6c5f3b0a789528694e, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h013c9a575382ff6881c908fb5184be7baf38edb0b06008592558efd57dd8fb9993c893800a6ac8c6d2e34ebfbeff43e63263f133868d0ac7a838f69aff26d60a3849, 528'h009d22ae7bca8a75a53214c3eece437fb28e05b076ec704d751a28a7ed7e529d5c5338be8c724afa547574a17f70510b2462748a53678e39752a688dc8cf39e886c2},
  '{340, 1'b1, 512'h0477828c9cc5710ded82ab21dfa5887f29edfb47548a5a99ff8315da76be5f67922c0a5de1cb7448a3a79b214889ffffffff7dc823ffb5d2fbcda33e63489df0, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01071ce5a19a09aacd43c7cacd58a439dcca4e85f94ea1d48a60f298ee01bb3eeb11d5daf545e7086486f8e4b518a15be69620ab920cf95c5c15ff178c903124fac3, 528'h01ad6eaeedece9a7592bd21508b2720f1b8c4bf55637b1e8a5ce5359775b980b21eb1d33e8ebf5c0b3d7829152a295b8a9a1343c25350e35f709936accc8ce08b0b1},
  '{341, 1'b1, 512'h17dfd1c9bfab4afc7d5ac126157041f4c4ca4a04aaf17c45e47857c384fb415e4362041ec3e91609325b7e4c9fb1a3ffffffff9d3efaa9406e392a0dea1ea309, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01bdae499160f4cc6cd163cf110bb1f9b421e8786a8ef9297e4b98fd508a1d14c50617c8d1a3de94fc8bd6c38055e4906b20fdcab6ef7bf9e7e5c98ef3e83e38ec3b, 528'h01ba867b8ee72bb7304ff83fc2d734749447420791d5609e0515de4e05fa70a83385a853cac6c47a075c8c61e4b65b9774574101cf4e081770f83ae1b7e727010ba3},
  '{342, 1'b1, 512'he2fc500440f25769bdfcc82cca36025aa6e5335d8653935dee2cc2a8e8a37c8a886885663c7da8224d2e807f62e1f039ffffffff2aa58c5c932713706022af2a, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0000269fc7ed89e554aa52b3875dc00bc140c1937d4f1b32e29da41ff241cdb9bd3058fc148f905982b8717b035e0db00ded7ebcb08572ec76bf0128411145d73091, 528'h01b4bd6bc4ba7befd5c305e018448a771b71fa1a11b3a2c6185dd6b8477c35eaeb4733fecd90f38ecba628f27c02f809191e993e1e7ff590383e2ec2afd08020b267},
  '{343, 1'b1, 512'ha5ce1cdebbed43dea085a592a1ef6c0881660e99434c6f3d6ec24874bb6cc9d56400958f7f95fdc15d3dcc870056263b85ffffffff9f3ace8f83061d0410f802, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01a5cecc0e572f5ee4eed6755d3230ec5a933c1fb0e35ae771a1fcf0dc880e1c159dd5b6d192dc377505048b7188de3feb815a81a4f30d9226cdc85f751dec1a0410, 528'h01ef4a743e1e16f0a60201cc1060625ede6f0936e7af90b42736281e89fe7f2de6aa3f25c68576da705d8b3f6d5d8a34d3073307ea198d1cc8d72a18ef25e90f31af},
  '{344, 1'b1, 512'h6ea638f8043673b9b6a79ff39b5d311774de5f4d697e5251ede52feecabba85d705f25c58b7c2efc844ce598d1428d22e4b3ffffffffc75b0ecb7283d80278f0, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01a92b43f57421e54d2528d305e7d5aac9a708e75a7d6fedb47908a4e3edcabdd836a2c4e8436f3b7b64895254536174d88c6dca143699522bc2dfdeebcbf38eb905, 528'h0093b0b99a89de72aca0c03e12724c2be323577a4629cb47fdda5b12b61ace0b9fdb97549d3d2a1dac15da66ba6389ee54cbc82c995b9f3aa3ae8474f4bb4b52da8a},
  '{345, 1'b1, 512'h7cd22c5fec3646707603f858ccd785676b3284b63652913e5581a60e0c262034285489fb945534b7f2578b3e64e7b956bb6586ffffffffc05edada940cffb928, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00a0400f255174ffb8548c29f5faa70e806bb6f6ca08a08753c85c5d145a555cc8e2df285af9985f2e729d4a99a734b7e7fc95560d546a067fda03529f56b2fe66bc, 528'h00d7fb60271d22ecb5d8ec904a9df1a416be706ce539e34650b8fc514d1dd7afebc1344c0c68c533c5b20ee249a77c075293b2d7efc8731c2e3619be59da871bb083},
  '{346, 1'b1, 512'hd289f68304c484efc5008425cbf00039a52c7b9d15476d36d58f1515d48a9ec94a850c121249365d7226fb6aad3a82c9eafe994affffffff58e8d36e4237022b, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h019207c7b645aa45c2722331f46e094f2eb0052075b8ac9414ad77baafd01d4d1fdc68344136fbce01edfa5627bfb8f3c128abb61072c74802192e89137c68d0cc31, 528'h00ff15b0218f81f0a848742f683cb4d1b7c517efdb8fcf8ac6a35e4971b35536851ed68de40a6e1a4a23bddb5b42efca23b91e91959a4f7e2afa196779c96c6c654c},
  '{347, 1'b1, 512'h792eae16afd3069393b20db2ed2e192ffd845b08e10d076d8eafc98744329d6279d31d55ad56a090712fe131358feb130a94bc4a2fffffffff97daeec1130838, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00aaf119702b9985354bbe3f6b6cda8c46151af4202546dfbe04d5f0ffd18ebe7b29d616f1c40376a412a52f4204b5a13e7f3e4304ead566fc41bf4b5fc0b84c8a2d, 528'h00d599deafd4fa2368cd072b854a3d53425d06adf3573e886b81248a7328a546ddc41caed38c6b1ffeaec9a98c940905cbffa87b936da980d4a9003da41e0c59c92f},
  '{348, 1'b1, 512'h51ae80a63d993770d8a5957111af53dabdf3abb9cf9908bc162ded716d3b3c5af2924c076e87c96249a4d7650253ff5112f8a2e7d2aaffffffff66e0e9175efa, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h006c09a59e71cf34f983f75dbb4724c4828a93021cee8fd7d92af6941ca8efc9c5ddda7c49a0e1777225782e09313e3091f056122e585c4eaa689fb2fdb1cb7848d8, 528'h019f0c5ff6b4638f4c33916db76f9d078bfa8f9e25ae00348e46bb32d777aa26155b82ea73a9e4e2f21f6a65c73ed6c6ab2101cef3524d45b9fc6ea1292f1986acad},
  '{349, 1'b1, 512'h100c883756f36d7c944d934c08932a99a1c2eb9892cc39a13a80b22aadc526ad755265f9ebbc8d0c1ccd31240299c71604332ff56592b7fffffffff1224308a3, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h014e791c42f3998458c5e17f895d25c85cb419195d65e5a0b9a42cf13ddd36959c73460f54aa840d2254355c6ac626f440cb3a84fba632262c9dc5cab31be7da106b, 528'h00abb97b682f01f45168403613a7e2ff82bb4a9fc20952a35d935428f71ddcc799c6d9085fe3230d72261d73cd082e8108523da7ba0b1691ad6ea63f5f4e8e8909f4},
  '{350, 1'b1, 512'hf4272253af2b51df321249280f3f3e62fb1e4a4a556f88bf3d5ae20ac5cc3e035e7b2141f9139b2f21d431068b8d5d96fcaad0f106289298ffffffff51777f01, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h013ded35ddff2f97780bbc60b8cec89855a35183a48f8fa6bbdc183994bf89021118cc019629df72112b2c529c023e7a5cfce253f7fdb49105d238680b64275a213c, 528'h009c92e7a0f71608e8d8cfab3f850f7fda1a1a1d056e72254469afe5ceec3c718e6a462e1346941eb08c105501647502c1a810a29df8b208da6a5b296b2bd1e98137},
  '{351, 1'b1, 512'h8bfa5531067a5cbc9bf002be2397bd10dd183d7ae47a02c0d0a7d87e1f94af93ea7365b711cfa611750ac963de0551c900dbad9cd8071b503afffffffffe6b6f, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h01d0d29756ebff02b71674fa4eae37557ccd51a036fb1eb0b7121b405e7fabd60592927d805b75815af1bca6e9d6c5484225bdd0ec7a40735da972fd5ff645d86f1d, 528'h008b9fe55357dc118070cf898973a64e7554b734e900c675541e20332a260ca51a23248d9b8f47ded811cfce556a06a71ba5dc5b873075f264a6843e675caf06a534},
  '{352, 1'b1, 512'h8a5409853b325b917b8a2aa1eb394767bb07fa82af11357e777f7404e0955bc9bb9cc5a918475c52df4772a1207e3ee4f3e3d3c8e68e84e10477ffffffffd35f, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h0165fb993f39d350ed60c8483dd6e4e6736591dea974ecd8ab027d3839b752322ee220d40bb6fc0b0d5a8c42928bde50f659b18f51f42fb2b1aa4583892a9114a0c3, 528'h00a8816c09d47138bf662da4ba25caf44e24185696d4914a7de2b2535f73b9afbd3ffa9cb0a86a115e4d9ac5be48cf7e8fe276466abdf17127bcc7aaf4d096008ca4},
  '{353, 1'b1, 512'h8e38a571ec826b9af00de0c523b6e073aaf9380cc64fbc86755f33f065361d8963ea2c42796ac7516f53d689e1da364bb7caf6b22a5fee81410646ffffffff7f, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h000b901c88ea699e715f6db864e23a676e7f7f2415ac1f850f2dde1ad0d3f9c92e8c5de66d45174d619955fae4b0dfebe49c583506481d28d30cbf58e2ac49f370c2, 528'h0144c97b688b9ecc07b84c68095267e17e48232922756609e9859d18d2eb7844ec925150c39f2b3a255c882be705e0a8e30e68e49fe7914dbcc3ccfbc1d467050f80},
  '{354, 1'b1, 512'h0f3ad12803aaf9bc615745a47da85dd90bff191d3e9441cc2cc96bf8c01f5e514b256685e3e48f01a98a5f27d20cd1c317a6f816ca8611fbc8891236ffffffff, 528'h005c6457ec088d532f482093965ae53ccd07e556ed59e2af945cd8c7a95c1c644f8a56a8a8a3cd77392ddd861e8a924dac99c69069093bd52a52fa6c56004a074508, 528'h007878d6d42e4b4dd1e9c0696cb3e19f63033c3db4e60d473259b3ebe079aaf0a986ee6177f8217a78c68b813f7e149a4e56fd9562c07fed3d895942d7d101cb83f6, 528'h00abbd9e77ef1e2a36c6b06f063d93effb8e852387a94bfdf8359b5c18708f90d9f4e9749fd45347f637546b08733789c988fda4f0309551bde813a0bb1a232adee1, 528'h0191165d58d153fec68f5cc83bcf5891e2e0ca9681204876e872453e9ebd45870b6878ee437e4d833c6ec54337b779acbf9f8202df510d269a710d0c43e4e07b040d},
  '{355, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00491cd6c5f93b7414d6d45cfe3d264bd077fc4427a4b0afede76cac537a7ca5ee2c44564258260f7691b81fdfecebfd03ba672277875c5b311ea920e74fb3978af5, 528'h0144a353a251b4297894161bae12d16a89c33b719f904cfccc277df78cea5379198642fd549df919904dc0cf3662eeab01ef11b8e3cb49b51b853d98f042600c0997, 528'h00000000000000000000000000000000000000000000000000000000000000000005ae79787c40d069948033feb708f65a2fc44a36477663b851449048e16ec79bf5, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386406},
  '{356, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00491cd6c5f93b7414d6d45cfe3d264bd077fc4427a4b0afede76cac537a7ca5ee2c44564258260f7691b81fdfecebfd03ba672277875c5b311ea920e74fb3978af5, 528'h0144a353a251b4297894161bae12d16a89c33b719f904cfccc277df78cea5379198642fd549df919904dc0cf3662eeab01ef11b8e3cb49b51b853d98f042600c0997, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386406},
  '{357, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h015f281dcdc976641ce024dca1eac8ddd7f949e3290d3b2de11c4873f3676a06ff9f704c24813bd8d63528b2e813f78b869ff38112527e79b383a3bd527badb929ff, 528'h01502e4cc7032d3ec35b0f8d05409438a86966d623f7a2f432bf712f76dc6345405dfcfcdc36d477831d38eec64ede7f4d39aa91bffcc56ec4241cb06735b2809fbe, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386407, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e91386406},
  '{358, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00336d5d08fe75c50946e6dddd36c550bb054d9925c8f254cfe1c3388f720b1d6500a90412b020b3db592b92ab9f68f1c693b8d1365371635e21bc43eaadf89e4e74, 528'h01d48d60319dfd06f935fc46488c229b611eecd038804ae9f681a078dde8ed8f8e20ad9504bcf3c24a0b566b1e85b2d3ed0a1273292ff5f87bae5b3c87857e67ed81, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe, 528'h0095e19fd2b755d603bf994562d9a11f63cf4eadecbdc0ecb5a394e54529e8da58a527bc6d85725043786362ab4de6cbc7d80e625ae0a98861aea1c7bf7109c91f66},
  '{359, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h006f8fadedbae63701072c287c633f9c0052ea1e6cd00a84342cc0f626210071576abfd0875664b0746cdaf2745effc18d94905b0fc9d2cad4ba375c0ea2298c8d1c, 528'h0150d128cb62a527ae6df3e92f1f280ea33248711ffe4b35c1b162a9508576860165e0ddc361d96fafcd2ff82776c743b9cd6845db61eb56739f5c4ef561e6c20d8c, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe, 528'h0015837645583a37a7a665f983c5e347f65dca47647aa80fd2498a791d44d9b2850a151a6e86fce7d7bb814e724ff11b9ef726bf36c6e7548c37f82a24902876ee19},
  '{360, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005e7eb6c4f481830abaad8a60ddb09891164ee418ea4cd2995062e227d33c229fb737bf330703097d6b3b69a3f09e79c9de0b402bf846dd26b5bb1191cff801355d, 528'h01789c9afda567e61de414437b0e93a17611e6e76853762bc0aff1e2bc9e46ce1285b931651d7129b85aef2c1fab1728e7eb4449b2956dec33e6cd7c9ba125c5cd9d, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{361, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00b420fb1fecdd9cc5ea7d7c7617e70538db32e6d7a0ad722c63580f1f6a1f5537eb50930b90fd6fdd9abd40015f746d2fd8adf945a75621407edb6863588e41979e, 528'h00295108a7e9d2191a287fd160bd24f498055dc9badbd61c6a89fede27b4f9d479d86a20b6dc07c90f008ebe68a0e0cc15a4a03b8cf990e4ff7ed6e3892b21c52153, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002},
  '{362, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0032b9a17c201aec34d29b8c2764e7c7f6aeef10fb61bf9837117fad879f8c6a22a300006d2018cf42b25898ffc9a1bf507352e59e6a52e627cda160e17ea2f46005, 528'h00317a89899b7cb3a0d33eafa02b0137a0fb1b05102b22b676f35b9ff6c050ddee9f185609ffb7f5165a769e440792b75044a43e838690d13f884aaae888bf5f86f0, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003},
  '{363, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0032b9a17c201aec34d29b8c2764e7c7f6aeef10fb61bf9837117fad879f8c6a22a300006d2018cf42b25898ffc9a1bf507352e59e6a52e627cda160e17ea2f46005, 528'h00317a89899b7cb3a0d33eafa02b0137a0fb1b05102b22b676f35b9ff6c050ddee9f185609ffb7f5165a769e440792b75044a43e838690d13f884aaae888bf5f86f0, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640a, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003},
  '{364, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0067dd456b52f82a5d4c4a71b3ea9302f62a852ddc04ad25b62fef1ddf657374fb4e80679ddf42d212f0711db32b626d8593bd70892e93ed0adb273157b6df187938, 528'h014d2c78509f3bd6f7d0fba4a90cb456286e267f5dd9d967842a6086884d66c7b2a932833470c721a4a728cd8486d15314232d801f17e3a6fd7068bdebacdf82c0b4, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e914b3a90},
  '{365, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0068d7b518214766ac734a7461d499352444377d50af42a1bbdb7f0032065ee6dc341ccf231af65250e7d13a80733abebff559891d4211d6c28cf952c9222303b53b, 528'h00a2f3d7e14d9d8fabe1939d664e4615c6e24f5490c815c7651ccf6cc65252f88bcfd3b07fbdbaa0ba00441e590ccbcea00658f388f22c42d8a6d0f781ae5bb4d78b, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100, 528'h01efdfbf7efdfbf7efdfbf7efdfbf7efdfbf7efdfbf7efdfbf7efdfbf7efdfbf7ef87b4de1fc92dd757639408a50bee10764e326fdd2fa308dfde3e5243fdf4ac5ac},
  '{366, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h011edc3b22b20f9a188b32b1e827d6e46b2ed61b9be6f4ada0b2c95835bee2738ec4dc5313831cce5f927210a7bc2f13abc02fa90e716fc1bd2f63c429a760ed2363, 528'h0118daad88fe9b9d66e66e71ce05d74137d277a9ca81c7d7aef1e74550890564103cc0d95d30f6205c9124829192e15d66fb1f4033032a42ba606e3edca6ec065c50, 528'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002d9b4d347952cd, 528'h0100508d073413de829275e76509fd81cff49adf4c80ed2ddd4a7937d1d918796878fec24cc46570982c3fb8f5e92ccdcb3e677f07e9bd0db0b84814be1c7949b0de},
  '{367, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h012f8b9863a1887eca6827ad4accc2ba607f8592e5be15d9692b697a4061fcc81560c8feb2ae3851d00e06df3e0091f1f1ca5ec64761f4f8bd6d0c2cab2a12102444, 528'h0174b4e34aec517a0d2ceb2fd152ed1736bc330efca5e6d530ea170802fb6af031425903fa6a378405be5e47d1e52f62f859f537df9c0f6a4a6479a0aadafe219821, 528'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001033e67e37b32b445580bf4eff, 528'h013cc33cc33cc33cc33cc33cc33cc33cc33cc33cc33cc33cc33cc33cc33cc33cc3393f632affd3eaa3c8fb64507bd5996497bd588fb9e3947c097ced7546b57c8998},
  '{368, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h008aed779a32b9bf56ea7ab46e4b914e55c65301cdbe9ea6e7ed44f7e978c0365989a19a5e48282fb1158f481c556505d66ff414a07003ebf82fca1698c33f2884c6, 528'h00a62426993ed5b177b6045e60b5fa1a1f8ce1ad5d70e7bc7b5af811dbf86e651f9ea02ec796ab991e1439bf07ffe2ac6052a8a0b0174d78a9441aaf4d8fc757d80f, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100, 528'h0086ecbf54ab59a4e195f0be1402edd8657bb94618fab50f2fe20fe5ebbc9ff0e491397ed313cc918d438eedb9b5ecb4d9dfa305303505baf25400ed8c20fc3fc47b},
  '{369, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0093697b0378312b38c31deae073f24a8163f086ac2116b7c37c99157cfae7970ab4201f5a7e06ec39eedbf7d87f3021ca439e3ff7c5988b84679937bab786dbe12e, 528'h01c6987c86077c05423ac281de6d23f6a685870e12855463770eccabc9f3a1d23cb2a0c15479420b5dd40fbdc9886c463b62ee23239df3a8b861c3291d28224f6057, 528'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000062522bbd3ecbe7c39e93e7c24, 528'h0086ecbf54ab59a4e195f0be1402edd8657bb94618fab50f2fe20fe5ebbc9ff0e491397ed313cc918d438eedb9b5ecb4d9dfa305303505baf25400ed8c20fc3fc47b},
  '{370, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h019a9f1b7b7f574a021fedd8679a4e998b48524854eefbaae4104a3973d693e02104fa119243256e3d986f8b4966c286ab8cb1f5267c0bbd6bc182aeb57493a5d5b6, 528'h0158b97eb74862fbca41763e8d3a7beb5fccd05565b75a3a43c2b38b96eb2ccff149c23ef1ac09fc455d808ff28081e985f9e172fc62d0900585172cfbff87383595, 528'h01fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138638a, 528'h015555555555555555555555555555555555555555555555555555555555555555518baf05027f750ef25532ab85fa066e8ad2793125b112da747cf524bf0b7aed5b},
  '{371, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01aa9f3a894b727d7a01b09c4f051b469d661de1e06915b599e211463319ac1b7ca8a6097f1be401d70a71d0b53655cdf9bef748d886e08ee7de2fa781e93ec41a26, 528'h01ba9ea67385e19894fc9cd4b0173ab215f7b96f23bc420665d46c75447bf200ae3ac7b42bd9b857fd1c85cce8ea9c8d2345e4687dd70df59f5149510735bb9c7b64, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{372, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01aa9f3a894b727d7a01b09c4f051b469d661de1e06915b599e211463319ac1b7ca8a6097f1be401d70a71d0b53655cdf9bef748d886e08ee7de2fa781e93ec41a26, 528'h01ba9ea67385e19894fc9cd4b0173ab215f7b96f23bc420665d46c75447bf200ae3ac7b42bd9b857fd1c85cce8ea9c8d2345e4687dd70df59f5149510735bb9c7b64, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{373, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h002a07f13f3e8df382145b7942fe6f91c12ff3064b314b4e3476bf3afbb982070f17f63b2de5fbe8c91a87ae632869facf17d5ce9d139b37ed557581bb9a7e4b8fa3, 528'h0024b904c5fc536ae53b323a7fd0b7b8e420302406ade84ea8a10ca7c5c934bad5489db6e3a8cc3064602cc83f309e9d247aae72afca08336bc8919e15f4be5ad77a, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd28c343c1df97cb35bfe600a47b84d2e81ddae4dc44ce23d75db7db8f489c3204, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad},
  '{374, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h004bb904073cb6da9e5028df54fc22cf5a9d5ca73a01feedd2b4ce43b87bfd4300a72bdf26b146b2e7b506c03c7a0ad4a7e3e67204dddca9b65d43560ffaf9bfd540, 528'h012b8895632e0406b78463fe1bc5360a3cf796fddda9db2b18ca9171558e6158fa4b0b1d0461d9a46b9b958d629bd62a29ee3942238e0fa83e932a66abb1b50c5f37, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd28c343c1df97cb35bfe600a47b84d2e81ddae4dc44ce23d75db7db8f489c3206, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd28c343c1df97cb35bfe600a47b84d2e81ddae4dc44ce23d75db7db8f489c3204},
  '{375, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h016454afca385eb53eaeaab711537d95c50e01268b100a22656adf5cedf68b4a78a6c14a70245df707f6565ce15948c2e38e3d90e05dda3188ab43a73f30dbc6bda8, 528'h0151dca6dc5aec84fa35c79f21365993f0b267ca486ea66c2186a52a3fb62b53501ce2822d4691fbc25cf27adb70734071be523b9231dd8d33a401dea00cf0ae30a1, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd28c343c1df97cb35bfe600a47b84d2e81ddae4dc44ce23d75db7db8f489c3206, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd28c343c1df97cb35bfe600a47b84d2e81ddae4dc44ce23d75db7db8f489c3205},
  '{376, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0060daf59638158ed9d3d7e8428501334764162f9be239e168fae9af348c30a7be1cfa4d9636c3bb621d7e0aa71446f8d4a37f2d43274a4255b226f612382f63152e, 528'h016e48300124a636b206fad4d0355862a852623799afee941e864d96dcbf55b801cabd6249b6f567506d5a503e7d03b4764c70fc44c5365f32c3603678476d62b09d, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad, 528'h000043f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc},
  '{377, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0051fe6a35a85070c7c29502a87672a38153d799aef734226b64d8fd3398621701117f0af9d9afaf6dbb8ca3007255dc79b0f41ed552512cb29207b15a01cdfdfaae, 528'h01a16c61277586356efadcb24764f21f574ef96f2caabc3f47fa66fb8719d7785824061c2d6d7a4bcb851540e62b2f00960b283eac7808d1813ef51b46e1149d3e4d, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad, 528'h01ffbc07ff041506dc73a75086a43252fb43b6327af3c6b2cc7d6acca94fdcdefd78dc0b56a22d16f2eec26ae0c1fb484d059300e80bd6b0472b3d1222ff5d08b03d},
  '{378, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00b4ffc0fff087607ad26c4b23d6d31ae5f904cc064e350f47131ce2784fbb359867988a559d4386752e56277bef34e26544dedda88cc20a3411fa98834eeae869ad, 528'h009d6e8ca99949b7b34fd06a789744ecac3356247317c4d7aa9296676dd623594f3684bc13064cab8d2db7edbca91f1c8beb542bc97978a3f31f3610a03f46a982d2, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad},
  '{379, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00809fba320fe96ded24611b72a2a5428fe46049ff080d6e0813ab7a35897018fe6418613abd860d1eb484959059a01af7d68cba69d1c52ea64ad0f28a18a41fc78a, 528'h01108acc5577e9e8962e2a7cea0bb37df1d0ca4050fb6cfeba41a7f868d988dbbcebc962986748fa485183f6b60f453ec8606f8c33d43767dddbbef8c412b2c37939, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad, 528'h015555555555555555555555555555555555555555555555555555555555555555518baf05027f750ef25532ab85fa066e8ad2793125b112da747cf524bf0b7aed5c},
  '{380, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0145130dca77d9674dfceffa851b4a2672e490e8fba8277622b0020e2fe9101e76933b0c01d248071f854e9bc523733936dc0b9930cbe154b9a402f681ee3c6cef6b, 528'h000d0c94b2ad28556643aa3d27523048d227a1de82f8a664707e75394d21da181bec82e1afb0e627539531affa849a2409bcac83fb786c351c88bac2fb2e4322e54a, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01556bfd55a94e530bd972e52873ef39ac3ec34481aebdc46680dc66723ab66056275d82bff85ad29ac694530bb2f89c36ce600ad1b49761854afc69ab741ce0294a},
  '{381, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00ed3e09809fe5985818f90592fd06e71d2c493d9a781714c9157cbafa5ba196b987fd49ae24274c76251c70b9f7970f1f713ad274590a702f463c73a0704831ce5d, 528'h00cac278297093bd9f9ac2d00bef3d67a01b43b28b9f829407264c738117438300c7704772976916ea102a776262ccf4222cc348c34aac683d8f00179a348323babd, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h00dcf9e7f441448a125b96d72b989d9f4dac7508c7e036f6080d4758e736f5e0636b0ff503f128a98d08e0ae189921065219d2cc3aa83e3c660ca0cb85e7c11a24d0},
  '{382, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h000ac2c5a4c79309a5132d5d7494befb3905d33fda5f80eeaf63775183aae7af108a3d97f3a441532cf6fac47f6c898329d69182e1fa07ce45997ebec3781c9ad741, 528'h0173a5b6b80a8b73d30ac97e1a4aacb773c1ad692c5ea63f68e373842782bd677864ff656cf8d1e6ec1e58e9a83856ef92677555916749fb95e800ae2e011618ca3a, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h0066eb57733c19a7003cf8253279fce41907bc4f127153c4576dd4814f8b335a0b51560b4447f0382c69b3fe509522c891f0eec3999ad2526835f33ae22a642843af},
  '{383, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01eb2a353dec6b460fbda49c67f431190fff6f195639c226ef8fefcbf191d72529a12cc5485b282a52704c1fd84529a1aa0ad794f96493e299718d2618a1b83a526c, 528'h01f704604d5b2b94a42bfc3ab93317d66a54de15258337433fc96a965d8e2d056fd1134b7989d7b3f709adc28227bdabc11fe2f359c6a6e5111ab43379ca25b66f2f, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h017106d1131b3300d7ffbc07ff041506dc73a75086a43252fb43b6327af3c6b2cc79527ac09f0a3f0a8aa38285585b6afceac5ff6692842232d106d15d4df1b66aa8},
  '{384, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01e43dfecc7e6caad03d17b407322c878f701c5add6eb2afcd786ff3803622dfbb6baa01246e1ea059f7b78842919b2507daa9e3434efa7e8d3ae6c35499f82d0ac8, 528'h018b0e4d6378222a07ccdb4214001f97b1a503d1aac3ab925ea64faa9c739ba04ee3480b147cb07f93edf40b6856a22f4159c3f5cd6c9e7165452907c8d02fab201e, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h006d1131b3300d7ffbc07ff041506dc73a75086a43252fb43b6327af3c6b2cc7d6ab94bf496f53ea229e7fe6b456088ea32f6e2b104f5112798bb59d46a0d468f838},
  '{385, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0141a4d714628c192b8ace1a42854da06e0e1ddb82a07618e4efb05d7095cd1eb65425078160594715eaf59fcb41c9e573fe10298c75c9e9135c775ca73f63d13aac, 528'h0089524b475170d4391cc032a0543ea22dab60ea07538f3a37607f0d4ed516634fde545e2f0a6ba8d0d2fe6aded0a771b4b134a5a280e54799fa476ef0ec87d44e1c, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h00da226366601afff780ffe082a0db8e74ea10d4864a5f6876c64f5e78d6598fad57297e92dea7d4453cffcd68ac111d465edc56209ea224f3176b3a8d41a8d1f070},
  '{386, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0147fbcc65d4818e029e0a3af13a1f7c90f0605a00cd0781200eb656a591d669a787620e6fc8cc594aa28a0b0f2939ec73472c494e09cecaf5f331dafd32d5ac31c3, 528'h0075432bdaeecaa0bec7feddc298c565723fb669ee76e38a4c5ff1701f1b38cda9dc9ac43bff18da2047e4dcd80c05a7bb7e7464829d608b68176b04c87f409f46d6, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h011b3300d7ffbc07ff041506dc73a75086a43252fb43b6327af3c6b2cc7d6acca94cb85df5e6c1125394fcd34f6521ffdaddd98f88a99fedcedd9384288bb793cf2f},
  '{387, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00b5b1c3998589b25c96a700bbd450d04da1f273df8053767a3b03ed1a763ed089c0de99bcf54d49c1520d3a09b845296f0445b3bd5b87918d3752cf651e0ff3007b, 528'h00e896380876b9419c56096914ff6eec01aee247eefef0741895f14ee280f360e11508c37826af82cd915b9002f046cb51008d9ead21124c591bd8265d1492b35ffb, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h0161be37ed5f748e06a89d72c4b7051cae809d9567848b1d8d7ed019221efb06ae81e1264ce49c5d29ee5fe22ccf70899002643aca7b99f57756f2639b6d459ae410},
  '{388, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01aadb41fadc35cf6d11a7c7d01d049b74b37677f04e1bd3dc08450fabae28adcd2d135f966616d283fb18a5e69eabfe7ec41e1a0edb3682f1d39f2af64a94d602b9, 528'h014ae81ebf5e3d2d0529479d4ae8eb05f4b42e519608466ad69e7662d6e9b236765f9be535c058f00f0866bbb4b172ef47a03cb97c58dde5750344bb293035f8e97e, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01e9bbbd64270b9668f7623ef7cbead5483eb07b883cf39fb6884aab67dac7958b0e03144357b9433e69adc696c86c63a23d35724cbd749b7c34f8e34232d21ea420},
  '{389, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01b706fc3f4aae5b86da261a66fbce47eb3b3e1e91544a40a9989fccf74154bbecac042dbbbf411a39090058b62c46fccd1d5eaba0c4879a688ea5fd0a7b4f9a0b4f, 528'h01eda01930c6b22745a97f2d59e182598dfdfbfdb463335293901de7fc9d49cf55ed7fcf5d767d4c22f89f171b4137c8415c3ed438089270c41f88eadef3018140e1, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h00924449b6c96f3758e3b085c079714f11f28d039b11699f0e9b3e7c553c8fc6c8f5212fec5eac3068713b8ec72fc6e2a90872b94e161a89822887f4a9bd5c9efd74},
  '{390, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0058a1fa96111bf30be76c3b8ba4435666677b6dd05031b5c4a840e1ea81f6025f70e1d395ef63cb59fa71e3674cb678f7250887f5d734e3ec377dbe3ae637d24f82, 528'h007a4eaf02cc57e658b5b9fa08ee30e0ef5b3429bb5a10438b0e05bacaebc60317010a334d7f896028aef620f5d9c7cabc38306e032b1b91c2376c3fef3e455a10df, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01554a01552b58d67a13468d6bc6086329e09e5dbf28a11dccbf91ccc6e2a4cfd4e6a2c5278791c6490835a27b6f7abb8a690bb060de3deb85093d3ae16482c84f64},
  '{391, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00303ba5ef90b05110002fdf74d2b8d4c7ab189c64004859c69d7c4730fcacb5f4d9b761ae987d1f3b63bb3ecb78aeecf4a04ff60f5f367a96ac2da8da27a3687a3e, 528'h006673d0d4ccd4c3ce1abc9980fd1885002c3e7b86078214caf7f0962fa51e116363032d7a1b93c92a4d62827549d5a33e4e6b9b6c2ab6ad9c2a15e410c5b1a846b2, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h00aa9402aa56b1acf4268d1ad78c10c653c13cbb7e51423b997f23998dc5499fa9d2f403c78b645cfba4eb78f595fe6d6f01dbaaf803f23ac263bf060baa74583abf},
  '{392, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00a94eea843a5c49637041598e30c381f7173bf8cd127f3caf5c16cbc728aa4d99173fb38d6a1b1ec21e40336e8d802249272b0ccbf4f8c3636ef66290a81b58fa5b, 528'h01116c23464fad61df8d2d5d1250a5a4c427e9c58e2cf1d059cdd88a7c34984fdd22a4cf18411e1b0224d444a5bd39d5fc97fc0b3648600f19d6ab80aa6a7c083a17, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01ffde03ff820a836e39d3a8435219297da1db193d79e359663eb56654a7ee6f7eb996c8ef12f62344ad211b71057928f96ae75b58e23026476cfc40ed0ef7208a23},
  '{393, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h014f71d2ca5bd2051336854657f09a1fab14c7f2f7865d71bd3fa354bf27b69dc8738972140553b525658b6fd203cc05ca0822e0904bad21b632e0de74a2ad3f0e72, 528'h004525f90519f9497425460b31cbb69ab3701a9ea68aaab72c6d65d364d0f0ed4d0524280f113bd69ef1ba9825202b10287a088c4bf30debecb720ac0739ec67434d, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h013375abb99e0cd3801e7c12993cfe720c83de278938a9e22bb6ea40a7c599ad05a5d3c8e5e5d7b3e16a99e528ef0ce91be0953cb1a9adf757f257554ca47ab053dc},
  '{394, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01d2ecad921dd100a8dc1a7b824b0ac6c9b654ab179833c2881ce237f1b8497ade851302cf50ea5ea169c2a50c0c09cb6ea539a7290a0f3437044b7a2e9ca8d40500, 528'h003fd5651535dcba1f331981c216a1c7d9842f65c5f38ca43dd71c41e19efcac384617656fd0afdd83c50c5e524e9b672b7aa8a66b289afa688e45ca6edb3477a8b0, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h005555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555554},
  '{395, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0165d67972a48fddc2f41c03f79ab5e0d42fd0992c013ead135c3394049645e26ad7c7be96510df59ba677dc94f1146e8e8e8fbe56debcb66920639581956b92b4d1, 528'h008aeb66ee0be18abaa909a973c70b5749d688f8e2cd2e6e1613af93d0033492d26a6e82cfb80ac6925ac6bc79b984f73e3ebbff2f223a38676891c1ecd784a8a789, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h009f57708fa97eba94c6d4782cdd4e33bb95c1353bde095232e3e2bab277bb5d2b48f55a53ffe928d034c29970a9e5f384a003907d3d9b82a86817cc61fb17f4c59e},
  '{396, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h018cd11252f0a434f446d3af18518c6b84cb0b7bf33758b4d83b97c2a56e0037b54d57d2b0b842e9c17d70504e01896389c066db8f2bfec025259a51dff514668308, 528'h01cca54365156c59e2c73c17664f09fcdcfd5b910f9ab48d0899b6a7064de8b80fc7a992e47ee7f23ec82fd80179a19f4cf89b4c02b7218f435298da5d322a982c1e, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h0068d98fa90736eff3e90f8fcfe50838b6fa0bf2cde77bc51e3f41019c8006f4e9cbaeadce7dbb44462da6425be9cfdaecb234c41749ce695be1b5ead2e6b1205f35},
  '{397, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01d6329a8afdea27cf1028a44d19c3c72927590d64628775f324514c81de301aa9be9c775c53a6349d1cbd5ecfc7bd39b373e613a10c1439441b141430fdadac168c, 528'h00071342d63dba901b93bdc444a1fe2ec6a15108bdf49eb1dfd218373884520d84bce03c5012f5837051cb8abf6a0be78dfdfeeb3a5872dff75b3f874faa6d2243bf, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h00e97ae66bcd4cae36fffffffffffffffffffffffffffffffffffffffffffffffffd68bc9726f02dbf8598a98b3e5077eff6f2491eb678ed040fb338c084a9ea8a4c},
  '{398, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01c963b64cdc3ecb1c35cda5ced9419ac146b060adb04c638cf6b66658013cb25e915a6ad0055668342881ed27f438b50ae4bb86ae3c7c02b727a130c77bad698008, 528'h00481bfffaead856b4137fd4268ecd74a6c2d4bd6cd13998ce7f0e828b220135d8df23253e681dc90673e0537e7590769a2a441aaaaa3a9901c4fbe44fa9513951ef, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01ae66bcd4cae36ffffffffffffffffffffffffffffffffffffffffffffffffffffb3954212f8bea578d93e685e5dba329811b2542bb398233e2944bceb19263325d},
  '{399, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h005dfbc867d53c57b2945502b8e56d96ca2d4d485aa33452200a2f4ba16042357976afeecf3e63b2fdcd5cdd76076c1a73e496caf9d6de3e8831d955d138e05884ae, 528'h01e04aa0b5360a0d3badd0120fbb8cc42a38bf1c61755d00858e40e4b10da4ea2575830dc92e312c20af2b8b167d7a58d178661d48cd932fe47a4bc7145e620ae22c, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h015ccd79a995c6dffffffffffffffffffffffffffffffffffffffffffffffffffffc2121badb58a518afa8010a82c03cad31fa94bbbde96820166d27e644938e00b1},
  '{400, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0078be6c43e366cf63ddc4235e8b969386e95012fbca5cebf1b0a6fe3c03c1257df7cf47b002eb6c4497f310bff6131b5ccb54fd0e8ee7fcf6b49d487e1b54508f68, 528'h009b61a547104c8516e0dc35d3d17659ca098d023b0593908fe979c29e62373738a3c30094ba47105a49edbc6e1d37cce317b49d2701470eeb53d9b24dce9d809166, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01cd4cae36fffffffffffffffffffffffffffffffffffffffffffffffffffffffffae18dcc11dff7526233d923a0b202cb29e713f22de8bb6ab0a12821c5abbe3f23},
  '{401, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0093f68961005f3040dc1a8ff1416c917bdcc77f1dfa85506c3bb62dac47f7be9529b4cbe57dd2c19e860bd2a0db71d47ef1eca8a20bfc3e0bc5e05c8303001c1960, 528'h002b9a3d45f2f5120fee06445f0d34e6138e3ac5b16d2a22f0460cea258c368ca9e478eb7b8253e7c6f2f7250fdc7dcd7243761f8d56f2350ac51e47ee063f41da31, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h0022e8ba2e8ba2e8ba2e8ba2e8ba2e8ba2e8ba2e8ba2e8ba2e8ba2e8ba2e8ba2e8b9c4c3f73cc816143fac3412b62de4c63db08f8c57e4c58c31f1b457ca5e57e20a},
  '{402, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h002d2d7d40bf17c4e8b18757e451ddded95e6b1007cd144809d21af31353b03038372c4af204d4414b71060b48b3a8439c632809bd33c4736263044405a1ad766e36, 528'h00bb0c5a8848f93fa3e85376b012bf064e303746529a673b852bb5a969c24c0156a8dd26242d0aad4bae43e23631b01fb9d050f9744b59f3b52b1c572217a1d70588, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h010590b21642c8590b21642c8590b21642c8590b21642c8590b21642c8590b2164298eb57e5aff9343597a542d3132f9e734fdc305125e0ec139c5f780ee8e8cb9c2},
  '{403, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h018ac11dfe62d1f2a8202732c79b423d29f43bec4db6080a220796a10f2685f92c71c7f72d9da0a8acb22680cca018eba2e8ba3bfde1db9a4ef3b97da16474364e96, 528'h005aad3b286707bd3ad07a060cabca49c53de4f56c05a0a8de40fd969d7d4f995f7c6701fe5c5321f85318b98be66251fa490088fd727da2454e00b3b94dc6e1241b, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01a4924924924924924924924924924924924924924924924924924924924924924445e10670ed0437c9db4125ac4175fbd70e9bd1799a85f44ca0a8e61a3354e808},
  '{404, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0051b2c3e0494564ed48ed3479b596ea4078240550a3c28da33d71d259e8e623e37ab43f396c49363f31c8de8a4644d37e94ed80e0dd4f92c3df2106e2795c2798b8, 528'h00a530d5e961f0696bbeb962aca8e71f65956ae04cdc22a4ac65146943e99a4a2fdb477df75aa069c8dd37a5daaea3848079a6a7bc03e0faa3d65d42f8053db2078b, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01d5555555555555555555555555555555555555555555555555555555555555554fa6dbdcd91484ebc0d521569e4c5efb25910b1f0ddef19d0410c50c73e68db95f},
  '{405, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01ba31a6f9c2d227da57de00759e2e844d607bc9bd92bcdf282006884dc347c9284f0dc0623af1e9db22117364a7a80a5b067efa19b204dac8faf2230d80b704addc, 528'h00d88b761cd3a4b0947bfc17e204b4d751f76880a82c9b7c6fd93ded55883c995002d8b8bfff1e021189c08d829d16b088f4fb39ad9456eafbc77c20353bc0f3c038, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa4fc31322e69da41162a76abf3a1b4507ae66074633446f259661a61c93be30eb5},
  '{406, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0137bbb48ef281133849ed723f5662a19fff9cc7389a0170d311bd34f4dbdc656246db695ea0712d8aceff9d1d0ef7921ec2e3f8b533e4ca122f9f7f446073889334, 528'h0163e4500d998095f60fa3fed4149d2d9b5b018e03eb5344efe8ffcc1c7d276e7401a4df639c4ab108820062495471be7b29398aadbae440a9bdcd55cf0bb5d96f79, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h017ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffa51868783bf2f966b7fcc0148f709a5d03bb5c9b8899c47aebb6fb71e9138640b},
  '{407, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00726dda8b7b6ed25f97f1fc6c3ccf554d60fc71e4fab2a578286d32612e7f3e669faed0b97619aef2d5aff9c8ffd987feddc0d6c38b7eec028191400874803f498b, 528'h00c0b8870c612e06c13c57ed6f7ef3d53b5e5fa2db62707b034b5ec13fb47018e31da7ecc991d575943468d701e118eca33122cf6d394b8a6ec0f45bc09701603a26, 528'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 528'h01346cc7d4839b77f9f487c7e7f2841c5b7d05f966f3bde28f1fa080ce40037a74e3001a2b00bd39ee4c93072e9963724941383cf0812c02d1c838ad4502a12c619f},
  '{408, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h016fce9f375bbd2968adaaf3575595129ef3e721c3b7c83d5a4a79f4b5dfbbdb1f66da7243e5120c5dbd7be1ca073e04b4cc58ca8ce2f34ff6a3d02a929bf2fc2797, 528'h0083f130792d6c45c8f2a67471e51246e2b8781465b8291cbda66d22719cd536bf801e0076030919d5701732ce7678bf472846ed0777937ed77caad74d05664614a2, 528'h0090c8d0d718cb9d8d81094e6d068fb13c16b4df8c77bac676dddfe3e68855bed06b9ba8d0f8a80edce03a9fac7da561e24b1cd22d459239a146695a671f81f73aaf, 528'h01150b0fe9f0dff27fa180cc9442c3bfc9e395232898607b110a51bcb1086cb9726e251a07c9557808df32460715950a3dc446ae4229b9ed59fe241b389aee3a6963},
  '{409, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h016fce9f375bbd2968adaaf3575595129ef3e721c3b7c83d5a4a79f4b5dfbbdb1f66da7243e5120c5dbd7be1ca073e04b4cc58ca8ce2f34ff6a3d02a929bf2fc2797, 528'h017c0ecf86d293ba370d598b8e1aedb91d4787eb9a47d6e3425992dd8e632ac9407fe1ff89fcf6e62a8fe8cd31898740b8d7b912f8886c8128835528b2fa99b9eb5d, 528'h0090c8d0d718cb9d8d81094e6d068fb13c16b4df8c77bac676dddfe3e68855bed06b9ba8d0f8a80edce03a9fac7da561e24b1cd22d459239a146695a671f81f73aaf, 528'h01150b0fe9f0dff27fa180cc9442c3bfc9e395232898607b110a51bcb1086cb9726e251a07c9557808df32460715950a3dc446ae4229b9ed59fe241b389aee3a6963},
  '{410, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0110fb89aff135edb801a1cb5bc49525b81dc74da45090d228122871814f489fdcb02ebee46b703e6b4e6af56c5024422b31fd4252c44d0bfd29d945de782d98543f, 528'h01ec425b4c4928e12b619227f1da6d0a9675070d9c5b49ca523050acb718e62643b0e5801543b76dc11f8d694ba09436d8391b477ad2c143ec50c2384c4f688512dc, 528'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad},
  '{411, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01c693a3fccbc9f625284239c2725f2a5c90b29b7ce3d07730f7de6031c9e74446d217888ae023aae23df6a4aa153f58c79597d57f42ce5c1354e5dc43a5eb311e13, 528'h015f99658443b2e39c3edcbcda70707fc5a4d39545eabe354816d09284a6265e47ebf0a47355828e818a767f8452a6d18451e0e3817a896ff404cb1611bfc4c4b4a3, 528'h020000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 528'h0066666666666666666666666666666666666666666666666666666666666666666543814e4d8ca31e157ff599db649b87900bf128581b85a7efbf1657d2e9d81401},
  '{412, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h017d7bf723678df574ce4366741e1d3787f834af9997b41c8260a074cb1f325d2bae9f8565dc6b51b6cb02dceeb5a1b774ee8dd7057c99e2d94c3c71299a9ce0f1b0, 528'h0162c65632fff88bdbb17ce2525ccac8df37c501ab0e6626e273fb6cf99000424344c0ac539c9fd6c4f3d28876b257c010d347a45bb010cc058443843a758328d491, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad, 528'h0066666666666666666666666666666666666666666666666666666666666666666543814e4d8ca31e157ff599db649b87900bf128581b85a7efbf1657d2e9d81401},
  '{413, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01e06db423a902e239b97340ab052534ead37e79412c675bf0eb823999e6b731040bff2b0e4fa64edf3962a328921ea5ae4e8f4079eab439e12f92335dfc4863c07f, 528'h007ee9f0ecb409cb133c0cd08b85e840b076f3d615e1ef1393b5222338b227d768003da5f3ba1f72f6654ca54ac11c2ba91a6cb5883d6d1a82304ad2b79de09215f3, 528'h00433c219024277e7e682fcb288148c282747403279b1ccc06352c6e5505d769be97b3b204da6ef55507aa104a3a35c5af41cf2fa364d60fd967f43e3933ba6d783d, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad},
  '{414, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h015053744d53811dbed8880f38d3a34578a7f1c172ec65bd8ad8183ba0ae10093416107f3c942742bde60719949b2c4f026f43582125c99ed48cbc7c5a051a5a7448, 528'h00b36d4c91a2b0367c566b2c12981ce0fdbc3beb983717403f69bf4264fc6182478af0b236ff120bcfca116924c552abef6663b6023be1986b70206d9bb89b5ed298, 528'h00433c219024277e7e682fcb288148c282747403279b1ccc06352c6e5505d769be97b3b204da6ef55507aa104a3a35c5af41cf2fa364d60fd967f43e3933ba6d783d, 528'h00492492492492492492492492492492492492492492492492492492492492492491795c5c808906cc587ff89278234a8566e3f565f5ca840a3d887dac7214bee9b8},
  '{415, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01fb2e26596cc80473917dd46b4a1d14bd9a1ca9769dd12bfac1bff17cdc282e74c73a801ec1be83edfe4bfe9813ec943ac151678f0a9a0bf27d9ef308177eb0400f, 528'h019e03a5da3da67e6b8d068dbdacf091b9d5efadaf63f4a7e9c6b6ed0a1c9a5d3cbc3e0244d481066018fba7674a2b59139a5656780563bb4618014f176752e177e0, 528'h00433c219024277e7e682fcb288148c282747403279b1ccc06352c6e5505d769be97b3b204da6ef55507aa104a3a35c5af41cf2fa364d60fd967f43e3933ba6d783d, 528'h019999999999999999999999999999999999999999999999999999999999999999950e053936328c7855ffd6676d926e1e402fc4a1606e169fbefc595f4ba7605007},
  '{416, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h008422cea9dcf8ae01f7a157888f018a40a66461d3566ec4a4dfc89ecb3c2404be734d329137d630387b012d033221857d5bfb290fa8027640b4063072a3e5b14c86, 528'h0025a219e724b81814901a677a8bee9b716b33b16a5b65f2272956a46b5e8683dc896984309ac79449657a1895c9f62bde99c7f5e24ed2defbc9f8dde35ebd0bddc1, 528'h00433c219024277e7e682fcb288148c282747403279b1ccc06352c6e5505d769be97b3b204da6ef55507aa104a3a35c5af41cf2fa364d60fd967f43e3933ba6d783d, 528'h0066666666666666666666666666666666666666666666666666666666666666666543814e4d8ca31e157ff599db649b87900bf128581b85a7efbf1657d2e9d81402},
  '{417, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01bc19cf4b94bcd34114ce83c5f1a7e048e2fc4fd457d57e39b3da29f4766acbaef1c10cb13c796a6fffb56d6a392e47b6c74522df7fa02754c33d95b1a9a3c92a15, 528'h00f5744c2bed308cb4f41b512e632cd01d270ef1a0d3f47ea780e73c6a6c9ea6a996faef4d282896c64fa50f5b04e204c56b504bc122ffba7aea4574d7d7ab6303c0, 528'h00433c219024277e7e682fcb288148c282747403279b1ccc06352c6e5505d769be97b3b204da6ef55507aa104a3a35c5af41cf2fa364d60fd967f43e3933ba6d783d, 528'h01b6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db68d82a2b033628ca12ffd36ed0d3bf206957c063c2bf183d7132f20aac7c797a51},
  '{418, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h017b0ebce08b09f21e30d15e0edd9fcdf24ab4831ec8a65a3d1e38f72b15f0115da6ed1885e42fcfae31c0914b71e9df2cd106adc039a82810a92924dd154dc05da3, 528'h00c614d1afc4f63de3803bb5490a34e1e2fab9eb78422b21d377fc0d7f991b938c22f4d7dd665f8dd21fadde43172a55f80d05cc4557b6663f9e7a3fe490d25c5531, 528'h00433c219024277e7e682fcb288148c282747403279b1ccc06352c6e5505d769be97b3b204da6ef55507aa104a3a35c5af41cf2fa364d60fd967f43e3933ba6d783d, 528'h000eb10e5ab95f2f26a40700b1300fb8c3c8d5384ffbecf1fdb9e11e67cb7fd6a7f503e6e25ac09bb88b6c3983df764d4d72bc2920e233f0f7974a234a21b00bb447},
  '{419, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0004c3ec8d7d23ce74be8b9c7c27be869c23bafc6874ebc44f47e107422ab1e75ed09bebd7cb1ec4626e442bcf512a25c5ddde26eb08ba37506461830cf9241cbe9c, 528'h0050a1bc08f4ba8da1d641ac3891823ab519facd4159768b1c0738f0e23450f374e4d6de55cceed95722be635c5dc0023a1498862f87bfe61d77e20e592cc20bb2ca, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa8c5d782813fba87792a9955c2fd033745693c9892d8896d3a3e7a925f85bd76ad},
  '{420, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00a7c8204f2864dcef089165c3914dcc2c0896075870ca0bc1ce37856f80f23815b0c8f2ec05145c421049e80ec1e7694f9f04174bbef21bc0972e559cf222de7e1a, 528'h01ff1108c28f01b703820e1c0187912962ab23109618dfcb0c062ccee339002222a3f7dd8dd21675b0e20908fe5855ea876d6a9e02c5f5b793d38fdf79fb83603ea9, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h00492492492492492492492492492492492492492492492492492492492492492491795c5c808906cc587ff89278234a8566e3f565f5ca840a3d887dac7214bee9b8},
  '{421, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01802fc79fc8e55bce50a581632b51d6eec04a3c74ac2bf4fae16ce6c7efef1701d69f9c00a91ad521d75ac7539d54bf464caeec871456103dc974354460898a19c6, 528'h00722fc1f528506618b1da9f8b2edbdbdaf7eec02e8fb9203d2b277735a1d867911b131f453f52ccc4ced05c3b1bc29e4d20f1e6d34979faa688ce8003f79d8e0c95, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h019999999999999999999999999999999999999999999999999999999999999999950e053936328c7855ffd6676d926e1e402fc4a1606e169fbefc595f4ba7605007},
  '{422, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h01beb0b4c2e494226404fca4ad505ebfed13d184b1572683215b16173c29a4475aede47f266e0c9c4143137d3e0001f9f0148b689286a7c64e229458b824ed765836, 528'h0130205169783ed9ada9f3a193027ae4e21829ad4a71d05d969605c04f3231dabab03beb2fab07dd8323d7132755734f4e6d1fb43fc8a63bfd244160c23efb6c1429, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h0066666666666666666666666666666666666666666666666666666666666666666543814e4d8ca31e157ff599db649b87900bf128581b85a7efbf1657d2e9d81402},
  '{423, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h0121e59aaf26b8301f4fcc3e0a563c4104ae00b47c55b8945ce749116fdf6761d768bd50ed431e2b51e646fe4fe7dc2985b6aefa7f9441ea11840d2ace2f34293cb1, 528'h000cf1e1a46d4d637216e28abd124cc641ae7a673445d573856bc2fec58d86e5ed63bc2a7f2049234e335a7bee95bb2724fb1480c97c38cd0d296cbcc113de3f135f, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h01b6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db68d82a2b033628ca12ffd36ed0d3bf206957c063c2bf183d7132f20aac7c797a51},
  '{424, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h008e859e66d1237fdc928a4b954954fef565d203a0731d065d9df41a4fd3812b1cc2487053ea19ce839d200845952f80d80698771d83ccc1fc7f236dbee4c76b2bb4, 528'h005a04b24c88cd40233fb43c59ea5cf2cb9510d16b1168bc126db64aaf9ab07a7453208fde079095966272bf03bc3312c9b9bab8c795ae375e8a0e8dd81c924e7c27, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h000eb10e5ab95f2f26a40700b1300fb8c3c8d5384ffbecf1fdb9e11e67cb7fd6a7f503e6e25ac09bb88b6c3983df764d4d72bc2920e233f0f7974a234a21b00bb447},
  '{425, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h011839296a789a3bc0045c8a5fb42c7d1bd998f54449579b446817afbd17273e662c97ee72995ef42640c550b9013fad0761353c7086a272c24088be94769fd16650, 528'h000043f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00492492492492492492492492492492492492492492492492492492492492492491795c5c808906cc587ff89278234a8566e3f565f5ca840a3d887dac7214bee9b8},
  '{426, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h011839296a789a3bc0045c8a5fb42c7d1bd998f54449579b446817afbd17273e662c97ee72995ef42640c550b9013fad0761353c7086a272c24088be94769fd16650, 528'h01ffbc07ff041506dc73a75086a43252fb43b6327af3c6b2cc7d6acca94fdcdefd78dc0b56a22d16f2eec26ae0c1fb484d059300e80bd6b0472b3d1222ff5d08b03d, 528'h00492492492492492492492492492492492492492492492492492492492492492491795c5c808906cc587ff89278234a8566e3f565f5ca840a3d887dac7214bee9b8},
  '{427, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h00e7c6d6958765c43ffba375a04bd382e426670abbb6a864bb97e85042e8d8c199d368118d66a10bd9bf3aaf46fec052f89ecac38f795d8d3dbf77416b89602e99af, 528'h000043f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00492492492492492492492492492492492492492492492492492492492492492491795c5c808906cc587ff89278234a8566e3f565f5ca840a3d887dac7214bee9b8},
  '{428, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h00c6858e06b70404e9cd9e3ecb662395b4429c648139053fb521f828af606b4d3dbaa14b5e77efe75928fe1dc127a2ffa8de3348b3c1856a429bf97e7e31c2e5bd66, 528'h00e7c6d6958765c43ffba375a04bd382e426670abbb6a864bb97e85042e8d8c199d368118d66a10bd9bf3aaf46fec052f89ecac38f795d8d3dbf77416b89602e99af, 528'h01ffbc07ff041506dc73a75086a43252fb43b6327af3c6b2cc7d6acca94fdcdefd78dc0b56a22d16f2eec26ae0c1fb484d059300e80bd6b0472b3d1222ff5d08b03d, 528'h00492492492492492492492492492492492492492492492492492492492492492491795c5c808906cc587ff89278234a8566e3f565f5ca840a3d887dac7214bee9b8},
  '{429, 1'b1, 512'hcf83e1357eefb8bdf1542850d66d8007d620e4050b5715dc83f4a921d36ce9ce47d0d13c5d85f2b0ff8318d2877eec2f63b931bd47417a81a538327af927da3e, 528'h012a908bfc5b70e17bdfae74294994808bf2a42dab59af8b0523a026d640a2a3d6d344520b62177e2cfa339ca42fb0883ec425904fbda2833a3b5b0a9a00811365d8, 528'h012333d532f8f8eb1a623c378a3694651192bbda833e3b8d7b8f90b2bfc9b045f8a55e1b6a5fe1512c400c4bc9c86fd7c699d642f5cee9bb827c8b0abc0da01cef1e, 528'h01625d6115092a8e2ee21b9f8a425aa73814dec8b2335e86150ab4229f5a3421d2e6256d632c7a4365a1ee01dd2a936921bbb4551a512d1d4b5a56c314e4a02534c5, 528'h01b792d23f2649862595451055777bda1b02dc6cc8fef23231e44b921b16155cd42257441d75a790371e91819f0a9b1fd0ebd02c90b5b774527746ed9bfe743dbe2f},
  '{430, 1'b1, 512'hdc5e71048a56da7aa1bf5fad1ae227446663488d8a531d490c4b5efa048ca4651acd9a196d9b13ee2a1c74ad440bdd88f6a34a02fbfadac2f7ce869e64486558, 528'h012a908bfc5b70e17bdfae74294994808bf2a42dab59af8b0523a026d640a2a3d6d344520b62177e2cfa339ca42fb0883ec425904fbda2833a3b5b0a9a00811365d8, 528'h012333d532f8f8eb1a623c378a3694651192bbda833e3b8d7b8f90b2bfc9b045f8a55e1b6a5fe1512c400c4bc9c86fd7c699d642f5cee9bb827c8b0abc0da01cef1e, 528'h005adc833cbc1d6141ced457bab2b01b0814054d7a28fa8bb2925d1e7525b7cf7d5c938a17abfb33426dcc05ce8d44db02f53a75ea04017dca51e1fbb14ce3311b14, 528'h005f69b2a6de129147a8437b79c72315d35173d88c2d6119085c90dae8ec05c55e067e7dfa4f681035e3dccab099291c0ecf4428332a9cb0736d16e79111ac76d766},
  '{431, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 528'h012a908bfc5b70e17bdfae74294994808bf2a42dab59af8b0523a026d640a2a3d6d344520b62177e2cfa339ca42fb0883ec425904fbda2833a3b5b0a9a00811365d8, 528'h012333d532f8f8eb1a623c378a3694651192bbda833e3b8d7b8f90b2bfc9b045f8a55e1b6a5fe1512c400c4bc9c86fd7c699d642f5cee9bb827c8b0abc0da01cef1e, 528'h014141e4d94a58c1e747cbd9ee6670a41eac3c26fb4db3248e45d583179076e6b19a8e2003657a108f91f9a103157edff9b37df2b436a77dc112927d907ac9ba2587, 528'h0108afa91b34bd904c680471e943af336fb90c5fb2b91401a58c9b1f467bf81af8049965dd8b45f12e152f4f7fd3780e3492f31ed2680d4777fbe655fe779ad897ab},
  '{432, 1'b1, 512'hd296b892b3a7964bd0cc882fc7c0be948b6bbd8eb1eff8c13942fcaabf1f38772dd56ba4d8ecd0b626ff5cef1cd045a1b0a76910396f3c7430b215a85950e9c3, 528'h012a908bfc5b70e17bdfae74294994808bf2a42dab59af8b0523a026d640a2a3d6d344520b62177e2cfa339ca42fb0883ec425904fbda2833a3b5b0a9a00811365d8, 528'h012333d532f8f8eb1a623c378a3694651192bbda833e3b8d7b8f90b2bfc9b045f8a55e1b6a5fe1512c400c4bc9c86fd7c699d642f5cee9bb827c8b0abc0da01cef1e, 528'h0008135d3f1ae9e26fba825643ed8a29d63d7843720e93566aa09db2bdf5aaa69afbcc0c51e5295c298f305ba7b870f0a85bb5699cdf40764aab59418f77c6ffb452, 528'h011d345256887fb351f5700961a7d47572e0d669056cb1d5619345c0c987f3331c2fe2c6df848a5c610422defd6212b64346161aa871ae55b1fe4add5f68836eb181},
  '{433, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00304b3d071ed1ef302391b566af8c9d1cb7afe9aabc141ac39ab39676c63e48c1b2c6451eb460e452bd573e1fb5f15b8e5f9c03f634d8db6897285064b3ce9bd98a, 528'h00000000009b98bfd33398c2cf8606fc0ae468b6d617ccb3e704af3b8506642a775d5b4da9d00209364a9f0a4ad77cbac604a015c97e6b5a18844a589a4f1c7d9625, 528'h011c9684af6dc52728410473c63053b01c358d67e81f8a1324ad711c60481a4a86dd3e75de20ca55ce7a9a39b1f82fd5da4fadf26a5bb8edd467af8825efe4746218, 528'h0034c058aba6488d6943e11e0d1348429449ea17ac5edf8bcaf654106b98b2ddf346c537b8a9a3f9b3174b77637d220ef5318dbbc33d0aac0fe2ddeda17b23cb2de6},
  '{434, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00304b3d071ed1ef302391b566af8c9d1cb7afe9aabc141ac39ab39676c63e48c1b2c6451eb460e452bd573e1fb5f15b8e5f9c03f634d8db6897285064b3ce9bd98a, 528'h00000000009b98bfd33398c2cf8606fc0ae468b6d617ccb3e704af3b8506642a775d5b4da9d00209364a9f0a4ad77cbac604a015c97e6b5a18844a589a4f1c7d9625, 528'h007c47a668625648cd8a31ac92174cf3d61041f7ad292588def6ed143b1ff9a288fd20cf36f58d4bfe4b2cd4a381d4da50c8eda5674f020449ae1d3dd77e44ed485e, 528'h01058e86b327d284e35bab49fc7c335417573f310afa9e1a53566e0fae516e099007965030f6f46b077116353f26cb466d1cf3f35300d744d2d8f883c8a31b43c20d},
  '{435, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00304b3d071ed1ef302391b566af8c9d1cb7afe9aabc141ac39ab39676c63e48c1b2c6451eb460e452bd573e1fb5f15b8e5f9c03f634d8db6897285064b3ce9bd98a, 528'h00000000009b98bfd33398c2cf8606fc0ae468b6d617ccb3e704af3b8506642a775d5b4da9d00209364a9f0a4ad77cbac604a015c97e6b5a18844a589a4f1c7d9625, 528'h01e4e9f3a7b800de63407b8703ac545226541c97a673566711f70e2b9ccb21a145ad4637825b023d1ea9f18e60897413711611a85c1179bff9c107368f1c1b61c24c, 528'h01de948ee577c3d4e4122a52ecccac59abb6fa937dfb3e4b988cb243efe98740309452ba013112b225b3b1b1384d5f68796845199a2602a8d4505a331b07d101188e},
  '{436, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00304b3d071ed1ef302391b566af8c9d1cb7afe9aabc141ac39ab39676c63e48c1b2c6451eb460e452bd573e1fb5f15b8e5f9c03f634d8db6897285064b3ce9bd98a, 528'h01ffffffff6467402ccc673d3079f903f51b974929e8334c18fb50c47af99bd588a2a4b2562ffdf6c9b560f5b528834539fb5fea368194a5e77bb5a765b0e38269da, 528'h00b6cf64861a2b16e33976095dbf45a592c7c24228c4a1dd727f303d5eeb87e5388ad05c328f824c40abd3e6ce003fef5cd59dee0069ad6348ea6e57f90f6bdc0a82, 528'h00228181c180366e5451dfef3593ce664804cb42d5a8d5046b816b3daf6602fafd9ac2dc24b8c93a10024480882558b6ad3d9e905923dcd0fd2a11964754a9b46b8f},
  '{437, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00304b3d071ed1ef302391b566af8c9d1cb7afe9aabc141ac39ab39676c63e48c1b2c6451eb460e452bd573e1fb5f15b8e5f9c03f634d8db6897285064b3ce9bd98a, 528'h01ffffffff6467402ccc673d3079f903f51b974929e8334c18fb50c47af99bd588a2a4b2562ffdf6c9b560f5b528834539fb5fea368194a5e77bb5a765b0e38269da, 528'h0093c8f766827d6dc15c810fa30433153a5e742859205ee8389fbf695c8840dc917440870acc5b160087ffd0cd9a6081029c60a7c26d5e8aa9a0570f4efdeb13dea2, 528'h012ec3bbf75a0ad3df40310266648a36db820217ed7fa94e9c8313e03293ef4f6a40e736fb8f208ad8fb883ca509d48046910523645459c27829d54431463b2548c7},
  '{438, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00304b3d071ed1ef302391b566af8c9d1cb7afe9aabc141ac39ab39676c63e48c1b2c6451eb460e452bd573e1fb5f15b8e5f9c03f634d8db6897285064b3ce9bd98a, 528'h01ffffffff6467402ccc673d3079f903f51b974929e8334c18fb50c47af99bd588a2a4b2562ffdf6c9b560f5b528834539fb5fea368194a5e77bb5a765b0e38269da, 528'h0152388c6da66164b706b41dd4dd48176d6eaf6525f876ef0ff2d147f6966ebfadf1767fa66d04203d3ec9c937a1f0c945aed953e34be444c219fd3b94d3277aa652, 528'h01658c1e5b2e563a49d11c883d05c491d628f0a92c3e3dc8db9a4c8d5f0dc846ac22af8b3c5fb5bbe2cfa98614dcffd87de1cee2c5912a5899505a0c5bcaa513e2c6},
  '{439, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h0000000002fba6a061201ea6b1ed4265163568735ebab78600cdf6a71101dc63beaf546d97a214fc6396793b014eb1aa7a728f53deb2ff9999a3808ddfed15e9629b, 528'h01993852dadc39299a5a45b6bd7c8dc8ec67e7adbb359fa8fa5d44977e15e2e5a9acf0c33645f3f2c68c526e07732fb35043719cfafc16063c8e58850a958436a4e5, 528'h010e89470f981d2c7c5c96587121a67323bb96ff2427739d0d885ea277293efa3b25c0bda04d81466198a3cbfc441f1b1b98f6bcdc2589d9d91a17a7899f70d0461e, 528'h017351b0da8c8d0e4aa0974669d190fa2f90aa50227160594dfb55755002365441de17ea42902128a6f81e554177ed509c0cec31fd5053fae03f62ff76579ba92bda},
  '{440, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h0000000002fba6a061201ea6b1ed4265163568735ebab78600cdf6a71101dc63beaf546d97a214fc6396793b014eb1aa7a728f53deb2ff9999a3808ddfed15e9629b, 528'h01993852dadc39299a5a45b6bd7c8dc8ec67e7adbb359fa8fa5d44977e15e2e5a9acf0c33645f3f2c68c526e07732fb35043719cfafc16063c8e58850a958436a4e5, 528'h011094ac23ca46a3e2b4ac3baae6504f1bfb3ddf2db9ab40eda32d8e0a05727998f8552a033bb05241e826a86a1d03014eae3aa5fe1a45caac1db3e8138b9cf59068, 528'h0147edb15a5080ee2f929f78b6ac86604aae51b674fa46eaae7fdfd90bf64d6189341155f4eba937eae74c9e480eb4fb7e6aafd4285e7fc503ee6ec20f0b1415be06},
  '{441, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h0000000002fba6a061201ea6b1ed4265163568735ebab78600cdf6a71101dc63beaf546d97a214fc6396793b014eb1aa7a728f53deb2ff9999a3808ddfed15e9629b, 528'h01993852dadc39299a5a45b6bd7c8dc8ec67e7adbb359fa8fa5d44977e15e2e5a9acf0c33645f3f2c68c526e07732fb35043719cfafc16063c8e58850a958436a4e5, 528'h01d876ae174da31e128babff9f1d15507660bdc7958750844dc4f4291f75a882a22f177f704be6067bf7ce8f06b8626d971e6ef5dcb666fa975c1e11126e04fccce2, 528'h01abb12630a68b669e6ad2d8d62654d75dfbc6b54a8e3a9c915be663e080ddcc348e57a10e2b1dd9f03e1b897796ad889b075e5919dc5bf37a112d92c693456e6457},
  '{442, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h01fffffffe1d5d52b31ca52f8947a35593edf164cd324f833b90935846c64db1454df9f028dc8bc36bb04cb7f0cceceba01a3844097f7c35eeaa81428db0cca63331, 528'h01b7c70277d0bf78a3c7b62c937f0cb2cad2565f5514f6205ceb1a193d4fdb45ba6e6cec07827bae0b16b8316c3539a15114d0de6d2de407fd7117551a70826eada6, 528'h004ed692af1ed1b4bd5cea3aa8ddc6f3f15d8a6ee0016fa0e8eb958580e7421832ecc0e387c34aafac6380bac419ea45c42ae6426af503847f22c49c2f456338c1a7, 528'h007aceadde02ace1668bc1a3360d34e125afde230f536c154d91e6c876bee1d34ae06edcbbca0c7cd17646840913164740b12e2e224fe3ef3dec6fd84a81b581c188},
  '{443, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h01fffffffe1d5d52b31ca52f8947a35593edf164cd324f833b90935846c64db1454df9f028dc8bc36bb04cb7f0cceceba01a3844097f7c35eeaa81428db0cca63331, 528'h01b7c70277d0bf78a3c7b62c937f0cb2cad2565f5514f6205ceb1a193d4fdb45ba6e6cec07827bae0b16b8316c3539a15114d0de6d2de407fd7117551a70826eada6, 528'h00e01094048fcf7a1e2ec66faedffc40f48c9c93514325bde6b4958d80f0413efde7eec1dc6de65f96009c069397e51da2eb1729efa287afd5552b25a9e427a6d836, 528'h01489e7e124f66942e642de992e60b3a86fcce576767719390c3a312fcdeaa560a7fbb0cabb35e05a6d6f3499160fd2dba12d29b613b16dec7494c950d65fdf11fa3},
  '{444, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h01fffffffe1d5d52b31ca52f8947a35593edf164cd324f833b90935846c64db1454df9f028dc8bc36bb04cb7f0cceceba01a3844097f7c35eeaa81428db0cca63331, 528'h01b7c70277d0bf78a3c7b62c937f0cb2cad2565f5514f6205ceb1a193d4fdb45ba6e6cec07827bae0b16b8316c3539a15114d0de6d2de407fd7117551a70826eada6, 528'h01d296292213380de133dc66eceb8bd857a5c468afe855c05da9db937373b51f9020ca11353415da76bb6af997a486d2370e31adcc0a4531952a3b59428678ee5943, 528'h015979a3c609c2c2099ae1b290da3d613b248e3a10de7ad770dffc82fb33e74fc3207533f97285cf4557a6407e9a775e59efeaee4264b2634933a6baf8c406f0c4a9},
  '{445, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00c7c8817bf2f0652a4a4b5140c773e261080a0a111395856e8a3350f5eb5612bd63b367b965e92e9538ea3b7908aef1ade4b68e17f9f9148495c167d1c4dd491349, 528'h0008bf0be2979abb8111fd0d768adcad774113a822c1bb60887053b5cf8c9563e76705a391ece154b5dfb114b20e351df4014bec19fa87720845801cf06b7fffffff, 528'h01ef8f785c51a25ae2cd93487b5c848d4af133217a91f51359c966e7538e68743578122df5830002f96f6fadb5bc44480e3b3b2c804e4c51cf95d059d5646c5cef21, 528'h01ba2276cc003e87bea37c3724e58a0ab885f56d09b8b5718f674f9c70f3b5ecfb4ad1f3417b420ec40810e08826efa7d8ad6ca7c6a7840348097f92b2de8d6e080b},
  '{446, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00c7c8817bf2f0652a4a4b5140c773e261080a0a111395856e8a3350f5eb5612bd63b367b965e92e9538ea3b7908aef1ade4b68e17f9f9148495c167d1c4dd491349, 528'h0008bf0be2979abb8111fd0d768adcad774113a822c1bb60887053b5cf8c9563e76705a391ece154b5dfb114b20e351df4014bec19fa87720845801cf06b7fffffff, 528'h0155978adc4b570d897511f5ecfb65a31947e6e989da17dea716625bb3fa7b92b853623eb0cd9ce2a5e2b4d8c1c2a90ec04fe79d012576ec728a45c5ce47c6d500c0, 528'h00f79fa8b94ee282a3d1815892cbf15d7ebdf62cb042c76bb3c710c23e32b75992cc249d84072198e4ed63d72435a07d2ed76f278d7399f61a5b5c997f45692fed22},
  '{447, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 528'h00c7c8817bf2f0652a4a4b5140c773e261080a0a111395856e8a3350f5eb5612bd63b367b965e92e9538ea3b7908aef1ade4b68e17f9f9148495c167d1c4dd491349, 528'h0008bf0be2979abb8111fd0d768adcad774113a822c1bb60887053b5cf8c9563e76705a391ece154b5dfb114b20e351df4014bec19fa87720845801cf06b7fffffff, 528'h01a2af29c58184ca861e7cd931f39cea064b199eee563f241cd5ecf6ebb2ade728f1be23cf007ebe8ef0c42d99f9f5190f6815446afc3043a820d7daf27e86b83b8a, 528'h01a2acd1822eb539383defff8769aad8bacd50cd24ca7aa6670671418110177808c3f4fbe6041b9cb898359ee61e04824adedd62b39fe5791907a20586333bd3c76d}
};
`endif // WYCHERPROOF_SECP521R1_SHA512_SV
