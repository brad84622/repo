`ifndef WYCHERPROOF_SECP224R1_SHA3512_SV
`define WYCHERPROOF_SECP224R1_SHA3512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp224r1_sha3512;

localparam int TEST_VECTORS_SECP224R1_SHA3512_NUM = 326;

ecdsa_vector_secp224r1_sha3512 test_vectors_secp224r1_sha3512 [] = '{
  '{1, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 224'h352507aabd0f9bc223e1ac97a4ccb33b9de8ad3df447037367aa413b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{2, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'hfba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{3, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 224'hcadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{4, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{94, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 248'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa52640000, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=248b(31B), s=232b(29B)
  '{95, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 248'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e9020000},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=248b(31B)
  '{99, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 248'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa52640500, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=248b(31B), s=232b(29B)
  '{100, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 248'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e9020500},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=248b(31B)
  '{115, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 0, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=0b(0B), s=232b(29B)
  '{116, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=0b(0B)
  '{119, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h02fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{120, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h02cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{121, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa52e4, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{122, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e982},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{123, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa52, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{124, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 224'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e9},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{125, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'hff00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=240b(30B), s=232b(29B)
  '{126, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 240'hff00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=240b(30B)
  '{129, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{130, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{131, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h01fba71f1257bc26e0a99d33024c3ffcddb31f81919d99d14a2a067ca1, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{132, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'hfba71f1257bc26e0a99d33024c41cf97f1ada11575df7ebf714e2827, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{133, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff0458e0eda843d91f5662ccfdb3bf19c52d996eac764357fb3255ad9c, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{134, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0458e0eda843d91f5662ccfdb3be30680e525eea8a2081408eb1d7d9, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{135, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hfe0458e0eda843d91f5662ccfdb3c003224ce07e6e62662eb5d5f9835f, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{136, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h01fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{137, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0458e0eda843d91f5662ccfdb3bf19c52d996eac764357fb3255ad9c, 232'h00cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{138, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h01cadaf85542f0643ddc1e53685b317a0a2389333e33734f17510e133f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{139, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 224'hcadaf85542f0643ddc1e53685b334cc4621752c20bb8fc8c9855bec5},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{140, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'hff352507aabd0f9bc223e1ac97a4cd9c98bd2fbcffe069da2e0b4e16fe},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{141, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'hfe352507aabd0f9bc223e1ac97a4ce85f5dc76ccc1cc8cb0e8aef1ecc1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{142, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 232'h01cadaf85542f0643ddc1e53685b32636742d043001f9625d1f4b1e902},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{143, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fba71f1257bc26e0a99d33024c40e63ad266915389bca804cdaa5264, 224'h352507aabd0f9bc223e1ac97a4cd9c98bd2fbcffe069da2e0b4e16fe},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{144, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{148, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{149, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{150, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{151, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{154, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{158, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{159, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{160, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{161, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{164, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{168, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{169, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{170, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{171, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{174, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{175, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{176, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{177, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{178, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{179, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{180, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{181, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{184, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{185, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{186, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{187, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{188, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{189, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{190, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{191, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{194, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{195, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{196, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{197, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{198, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{199, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{200, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{201, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{204, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{205, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{206, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{207, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{208, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{209, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{210, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{211, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{214, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{215, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{216, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{217, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{218, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{219, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{220, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{221, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{230, 1'b1, 512'hd5c6e3fadab991245367e0cd559cd915823b5bbc764608b2f8ac52e64f75e93475682903430b5f85d1ecf507e90a7cdfbd62318d36e44b64c2201df079778ed6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 232'h0091589658ccb7ceaf1f017492450e2915bb8d863bb7f398c8f5bc1387},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{231, 1'b1, 512'h0000000097ae34ada66084471ced074cb11f6012595501e4f88b5ab4526808fbaabfff3975c6cf53455cee950965a5b5b71310c8a1822cb5d15b513b43dc5720, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5ee27f9264ab53661d3a7b8c858300c6ee5978a30ae9b7e413dd680d, 232'h00f9e6c2aab2afed523b0172ba110b5b0d663a8f77220bb865cef20f4f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{232, 1'b1, 512'h4a00000000d34b9c928306129f1a8059b199049f30ffd4d5b9747c848b197497634fb5190298af2f6a90d273164d68431c984e0fcd3a810ccd7b95b5e0dcd21f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1bb6ce51b7e504ccd69a910a11a9c29ba77100d5bccb179de19a93dd, 224'h770a160b2635bb293c73a07fb1fd5e0314b50127ab3e70d1ab974de6},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{233, 1'b1, 512'hf25200000000600b35bfa47958845baa9428119e3a1641db59a3b72db0b47470dc44921ca1826d81bc2e78142986441cb6a6c15880383e1ed77282f966ad17de, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fd8a1f6ba87941c7a4cb8e9844fdba099bc30036cab0b82dce6802ac, 232'h009732c1f24fe6c3fa8113b756c6b7e1523375dbda788895018ebf0245},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{234, 1'b1, 512'h9e93cb0000000075ad177fa53827e2d0b2d93ab1e6b099c341864034009c13d5ae494352e6106d44bfde1e40f82fe0bc542154fd54365234bd13e0a0e4cbbf31, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00cfd828e8c9b0b17363136530af0a54a21a6cbffa7a20a257385118ff, 224'h7bc8791627fbb74a63a76c99f8bee1325987d0ab2a15b0d57604149f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{235, 1'b1, 512'h6d22e20c000000000726c9469eebfd2e764c9b4750557869e51bef687b0b07862ad496e4c6a056d46f5d244f5f10ad0005ded39047ab8247ec969c4e42ec2219, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h35e45149bdcdb55ae37a3a2937d2d03a65754e29605dcc5076d20aa7, 232'h00ba6f5eb05da4fa57217efcc03e8f59a35afb6c2043da8ffcdbfea1c5},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{236, 1'b1, 512'h5a5af3265a0000000025640fd363bfd88cc171f1966b1906138185d763f0ee7065ebd2a5813b79d02ca118763c60dcbda580f5ec322cdfb2c0a407e223f6b16d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3f5dfba448339287d1bac93830c83222408a7b511aad1d5f530dc6ee, 232'h00f4726edab91264106792e45f30c8b489d268291d3c2a166555dedfd3},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{237, 1'b1, 512'h6c0f86f08b1e0000000069a0652407ab389f7f275bee385294bfc2a7a9119905f5ce4e1af41b3850d665c942f16914cf903717ff47c4e186c7fc97496a068b91, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ab65412c5db588242b51644dfe78d72570e66ff846feb28112d2651a, 232'h0087ba5d4a58ed7999f502b79626b45a0fb19fd8e4572bc1b5d49b3b76},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{238, 1'b1, 512'h5ab9d448ee67ff00000000baa93e38832a2709f7238f9bceb67b53fea917f665de9153c44b7280e1a5674dee745f5350bb3f2259ea084b398cff74d33bded951, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009ee1f0edcf13e952d21c30fc3c0c05a7b7460603893d9530d8e90258, 224'h48efc43fc23f36f84970c9df74fb1a3e163e95a1063fb3ba966e3e8e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{239, 1'b1, 512'ha1eaba175145939e000000007804c10bafa1416c6dc9d3311f844fe42868c6bdf283b946814df78822f198d26d886ed4713421a20dddcd82a21333d922eb39a2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b279452ae24eb13cdf7f0854409a7a6c556ae42f590ad5eeb874e256, 224'h2cc96e8ff6e523c2f109080351c8e1542fe405227ff7542f2f924e95},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{240, 1'b1, 512'hb1fe8fe86f9994808c00000000f313a999ae7b5281bcacf933f05e4c8d526e761afa3141e9efefe959438620220c28bbad7047a6c1a98f95520baeb1d7af6278, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h398b59d0b6a7171d3518d1d3ef6796f10a14251aca5630fa32655741, 224'h4259d0edc9c2aabc09c37a69444df24a5191e21d387b98b080745279},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{241, 1'b1, 512'hfa3ef856182ec646db7300000000241a0e98fb88ce661de43bfd86f1c929391ee9ce6c05612b1609d6b8466a9c4d0af24ccb440f463cd18addf4674adb2f94ea, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c0604841fb5caf4f4f2f91fc7804729349f796adeb304486ea579e02, 232'h00dab85b543047ef1f2c2bf9feab25a6c1bfc89e5734edd69a3f8b09fb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{242, 1'b1, 512'hed19e69c6f4de76b35ce6c00000000ad94175b8ad5f1fb69995d7d87abd893772b81ff83fd6caa25d1fe69b0317ec4068cdddac49512e6bf12d9cd8ce9a951c7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7f5127a83c76554fe4fcc00ea6e62b14c8a675168e60ea9d6b1f034d, 224'h7ab4aca6a9315c795936fb41bcf46a4840a1e41a874ddb1ad5b550a7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{243, 1'b1, 512'h2e2e984df4c5b45f7e337184000000000600f130d66940e8b4c0c1030e71fb8df7efce69100b9174baac3e7c474054e875f26cc182e925a17f55688964033e9b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00aca0bf2ba598af7c37adb7617da4b1b2ef93b82b58f1161db8949ce2, 232'h0086d0e4743c15c74b1ab334e236fcf23976c731491c808cc55027521f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{244, 1'b1, 512'ha8f658c6632e4f474a6f1af1b9000000000048ac2a6121c8add714fb8cce854dbf1871b07a75008a42baa6cef01b4875eba4bc9327b41503cb36ac20f9354238, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5fd0efe2e36041cd23431bb85e2bc038994a706fb9a40ee8eaf1e664, 232'h00c494185ab2c6dff620f3d48bca6130d4d507e35a0090eb27f167bdaf},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{245, 1'b1, 512'he89af705f005a4e1c5983824150000000094795c26507ca965c1eaf5782dd829a5fb5464eae46688a19ca7fe5851291f76fcd7f7226131d74cb4dde6063215e8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0f173d33840439b0072b8315e735f3732a5657334b9d8a90faba6919, 232'h009be335cd9d18cf81a4faae6110f2532881ab57ec71ded448390ea224},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{246, 1'b1, 512'h9490ebaece67e31eca85b20871120000000077b2785e29958e0ab90faf8fcca953b142d51892ae5362246dc07a066ff6a4c9fed90a79fb59abdb7c8a888a9652, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h601f7bf10bf200a48369d222d9e4076671339aa98955de31ae7f4503, 232'h00a11b5f8b770d78aab8ce1918a60b496e3775e9f9097bdbc598c9e99b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{247, 1'b1, 512'hdf22c290212fe9b66a9c65575e7be8000000002b9d4a3251cc7b64eeee3e76b7e65ac253a2e3d18658634eacb7494688a1616feaa0bf8a6cc0edbdeaa4533490, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h07c32dca0c28e0b3a142944b4f37a1b9293175fbb577ce38642154cc, 232'h00e48d47870afc0f169327cfbacf49df87bf20a13f5c2a57854d214023},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{248, 1'b1, 512'hca6a7cd52432b20d8cc73c4e810dc325000000006ee638ed6bda85ccdf3b4606a300f2439910d382aa47f8e5839698e4bfa1756c5e93b3d6aee97edbc8ae7794, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ca328dba129ae9a7b273fd1b67d843e02d5bd2c4d77514891f2c08d5, 224'h44ae98af8fa9d515995ee5a6fdf56856c67c4fe5f8832781704dacfd},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{249, 1'b1, 512'hd912418a7d72e83ab66eed185bd627c70b00000000a88db442365b3ec21269abd09b4b2e040304518850835236add11fecca5a2c529f8bc4c06174a03b997830, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b00ebcedc8c30521024d15dfa14304f8c594ab8a17eb3df68393b2e, 224'h3a53183103dd1b1ef8631e7cafe510eac9ab4c10164df208c598e20f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{250, 1'b1, 512'hd8cdcf759b329e28b173d8582d7a91bb2d12000000001faab0678de44c1caaf5247d111c9e465596a89073d5492cadb0bc766620952c817f31a391f32fb27346, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4cf261aa6616509319653090abd707202026733fd64ddb14f2ab26d3, 232'h00d8e37fac62420a7e9944e4b319d5e73d03b87a589971fed7012ada54},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{251, 1'b1, 512'h91f07f1a3d4b600628f1754ae5ec28d43554a40000000051e8c4594c5a2e68bf2f497bfbc7e703e1b18398a0b5515a38d60284b1a2dfad8c9132a7b9a98db6eb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h504f2f50ca931e2a4f8cda0f08c2b79ef051677d76a08f1806c53af5, 224'h736248501f062b14bd3fee6528700d1a64a8ae30d7c76e1a92b66bad},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{252, 1'b1, 512'hc6208a5a5c6b71a957477d8c39b01e072a65ac1b000000005c6ec3ddb8ce20911bba1864112d3407082c700820f8676037efb40be95619c9f686163a4d0cdc5e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h79a548e4da3b3df4df774e7fb9dc4af0706635c454e9e23c2aa29752, 232'h00b74069eccaefba00a71f33b43f69eaa321dc58436ebafbcd574660b0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{253, 1'b1, 512'h7da7793b2bed3ce23ef7f1c04376791fa03f741f650000000008744fe10ac37fab4edf76492a339fe79e56ef75aee6c3169a0a61e3cb27e74666a4fe4184526c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h32377296ba47114b5f3dcff841416bca3e5e98d64dd987badc457655, 224'h29a37a143b47b029e256c7506a679ee8f1962ccbbb1c83f4088501b2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{254, 1'b1, 512'h48cd33f55583315ab2131d5db1f9cfcb0590b13a266700000000c9bd5d6fbcdf457e3bffd7b4875145a47be68b99a201b93b8685e80d61ce692a913be1183569, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h75d62c172f26e6e6831c233b49895c1a87c1ee3ef57b711856199e46, 224'h27830a8d1fc44993990a9d1b2b147ff8792b0b0823bc30fb012ce9ee},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{255, 1'b1, 512'h1acaa001f6ed1b1a5b0bbde85513fe0b7aed266bd9da3100000000dc1113ab87ae3bf815157a1926b7bc3f659934702113570c26bf1bcdf1c8492f79614e844c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fab62ad526e88f6b9ca7e2d23f38d9fcf861cb7cc275faa25ca6a09b, 224'h29b371dda6ef29f037181b9c3bd92c78578b43dddb74a029bea7f238},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{256, 1'b1, 512'hc6244ad67598a847488d31d513fc9dbd21d96307c296a4170000000012f527d2192eacdb6045c48c250e317b7fc62ea79321783ae0f400ea4a60b48c2a2fc495, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00939e3d378767fc069ee193f001f9c84e4f82dd40747e037df3fb200d, 224'h7db50ec017098cab3ad054530cee5238b0a315cdc80a3d8a7dd0991f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{257, 1'b1, 512'h90f9b7739bb1699b90bfdf7cef079649e3f08242a08d05026100000000d3a4568eccd5ef4d94de4885986b68670617f552b9cb2a6eed337392b49ad4d04a9dad, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1a71aa363800731f4c5a9f0a4235198a7658f1b425972ecac9a2a340, 224'h21b61939e575b1a5ff487473ba3803683c8b20e89844a55785630f89},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{258, 1'b1, 512'ha7ee711aed6f375a8a15680f30deb6946501624b70b47c79d5a500000000ee6f7f0f2b69cde1a389e3abe86e51efe844c8e4ee7c3b2a15925d8c9b8b296ccc53, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e7bd4ddedd412bdc8482f08e2df540576b1bf768933e1adda30ab963, 232'h00b7d647170f0cfb0324f9ec2e299403dc6cf1589be3dfc6fc228234f1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{259, 1'b1, 512'h9583a32b620d5614a1c36e06ee45750fd69ef561faeecded2ff5b4000000007bb68b2b419fd574ffe1760fa0203fb1718c4e5d8a798563fdd98439f37a56dab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ac96c0158f3f939d14238f744c9c2b5736c026db414c5d9c019d0562, 232'h00a27c8a34065c71b92af11d77dad533f9cc62667ea09d50057fbea9b2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{260, 1'b1, 512'hb6e404060dcf7182366941e77a0f0b43737232bbf9f73865863c271800000000a4ea51e31a92eede7497562eb5eff19b08310fdcd46cf3c22e069110aedc21a2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c526a888a4f74f01f037b7556955dfcae72266e5df55ac6cecbfb85d, 232'h00d85a5bc24cb73aba3188098c11f7087a39e5e62271e016cbca2b5588},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{261, 1'b1, 512'h57003aeb6ad8b84b54cdddb9243c65d8fd07ad1ffdd35f11c319f06394000000000aa9393490e8dcaf1c1e53ab5a7b2dfc0bd1dff4d0fc1e0c9dd5cbb035748e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h37206ede6a2f6bf468a91152503eb90837456a3b1d6c937b0efbf60d, 232'h0096d35182fd97438e4a978c2223eac6a4f7005926e895ff17d667a2da},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{262, 1'b1, 512'hb47f61cf42394fa1c4c8cea80b83e366e30a938140f793851af87bd3782900000000d7a39fae605c98c96e0a5b0e8a58e47c3b50d4905171c884a64239fdd901, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c42106cf72c3632d1d4f15a08b7bb72c57ae82c099953d324149b03c, 232'h00fad8d9d9da94259b719ff6b6c8e6ab24bb365602ec2ffe12fe0e02ec},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{263, 1'b1, 512'hdfe80a6b887fa09cbdc8bb94300a4ad38f0380331a18c0a0b62708e590dd3800000000d364091041bb72f35391e792802f5c23fd676d0775e56ac2e41880d92d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0fc1582e0b3ebe74b1fa4425e321a5b2d16b1c3ab060e98cf530defa, 224'h115eae025fa3422621a49fd78486ca245894a2d83c644e31abe21b5b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{264, 1'b1, 512'h16d0d407630fbd8dd9af18abdbdb902051c86b156254ecde6a5f0a5a1510f99400000000c202a44b1c172e1436f2252d80f9ab44794b22086f877c3bd4aa5fb3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c96588e99831484962138ee5cd487ddee8c2850c6e82db35f8d5ad4b, 224'h26ee8a0787b6c5bad7598e5d41e59880b32cfa125c8930fdb0c16480},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{265, 1'b1, 512'h519e4709f22b7ec44e321f4d403bdde7f532392786df003ecda243880f79f899f7000000000e3e6d749c0a602d959e0fd13a8a491554d233b9dcce6cac4ff3fa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d144ba07fe4c7f96353dc8b171384b4492cebe74c86cdffe6213f796, 232'h00c19fba0a58850f2ddad8ac81b404ef18f5b1b48198e48d069dd9c2ae},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{266, 1'b1, 512'h00ac9e66bf4db08b47a08e0b34e95e7ec2da8a82091479dabd2d57199b450dda70f8000000005b979f8077a5a74eaafe42ec70504f2bf8cd07aa23ef52c0321d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h48f0d2b55006514280ce7ad28336ab31a0536deef767f00ea3419b97, 232'h00918326b9337f76f3b3b3b789031e5c6d3000f7215b5d8eb38546797f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{267, 1'b1, 512'h2cd7eb20ee13fc351891dc4acccbc978161cc1b1e0cb95127485ff132176a972377cdb00000000add5eee3b407ef394da0255f21b9b8ca144d7e76fb075c6bc1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h44d3a182c9a8a207a5dcc2811e30eb26037bb5627870a1e3a754a1ef, 232'h0082a5978d2fdea3875cfea57b3178742c42ceedd3b396d5014185317e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{268, 1'b1, 512'hca402f2de7f990c5e1deee30d418810cd3a8707888fa5d54d3a5a0b3bab20144dbf37f52000000002a1f22f563f07cc9d066dfa8881777cdaf8a1ae4d43d6341, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00eeddc59d60f2757081c3b915984e739ce31ccbf184fef27d1025c711, 224'h686f704834047ae4b8beef8fcb67c94a05b7f4769d6dc98021c21d6e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{269, 1'b1, 512'h4386a89b56a955feed663fb88786a1c3916e8c65775648439638f2278c7d32c6d67f942e7d00000000d3a5ae2110db187684130f7aed62cb05159f8bb6eb1b26, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ba4c612540922f0a1b770d9373c518993fd445105057cf26c0aeff8c, 224'h4d6565ff7317d861b2f3c07df628a48d42d21a0ea99e8945486ca37d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{270, 1'b1, 512'h9a76ece71e15ffca113598c14654fea437156151bf5c8d47e15a6279ff965eedbe79fd4437f300000000148cc8ba720cd12a6cafa72448ec2cd6ad2852b2f703, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e67640a782681968972376b0fd72e54206af328a59be671e6158448a, 232'h00f2a76ed2674b1f9142f54c8fe76cb8dbff71f4df3775a2abeb120a2f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{271, 1'b1, 512'h24abce8b935764d6a61bf597db6c773145d5992485866070fe22cd0f6f871d53e72f6abbcac6ee00000000840dc44c1955185bfcf393a1786b04625904f03e85, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c520faa7574e13bec8b3f997ee9b844b6367d61d26ca84dfe4eb245b, 232'h00820be3e48aa4e569dd6d7a50e74d65b59fe603c9651dd3abe8ce9720},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{272, 1'b1, 512'h3fa9e7c5fd635a7b587b56e19e8921e7cdc6d8f6b1ff03b579b907ccc2dba540c1782d5c35e3aeeb00000000a610ad03b540240313bbf54453b27d3794341d59, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d86d566ff5fcccf3a356786e614b9340c242648c15ec4b670ea11f07, 232'h00abb0e7da14332b7742636b66b8b7beb2ac4a155fe6308aae6c70660b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{273, 1'b1, 512'h4025a46ad55fab109832d892d397d6e50c9c0aaf7136c275c259a6a61333a7e139b394a288148e32c200000000a3d26314f0694c5db5058ee34dfdd8fc2af9f2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6612d845fa2d59be90a0cd7f75a3509430ac8078317d385fbef568a5, 232'h00c5df1cd8920cd3b872e2335522bef8295cb544082d269b83aff84eca},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{274, 1'b1, 512'h1e2fbff1179de8374cc3b5f47b00ade36b6494b8941aa810476c8b40e3ad3d7f5f60d8ff0d13bdc7683d000000005b2a7c0d9bb60d8af2267c656e800069cee8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h098f5293e6122fd450e1f3182e6f2323b5878b39afa4184883977c3d, 232'h00936a9af99a3c54e1b94a04fef86cc7a16526fea66f6a1c3d40da1604},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{275, 1'b1, 512'h1efc0d2c8682584f2504efc8fb5fd2848583ab11c97a1ad1d23db89d7d853316fd159eb4e2cee6ee4f2eae000000003ec9bbec801c26e55e61dbd6364bed8027, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f5a524acbbade6852c29132c32d61b06707a388cb3cebd8eeb59d1ad, 232'h00d7de65c50b21a84e6f49b71fdaf977e3d2ee8fec008e477428b0857b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{276, 1'b1, 512'he68fbb72e90ec509836476f39f26d3f65c5deffafd5b86448457438ee0c621fc8f97e83c77ecd131ff1e33e6000000007c2a942574c7da923726d5304e0de79f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d7c5da509bf42983f7ef6d7578eb297f58b51b2c47001c6fdf3aafe8, 232'h00c6ac0690050f22e9fb9f0fdaa24bd1558f793a0a9a5692f8e57959fa},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{277, 1'b1, 512'h90bc23f7e48f29ee5cf5bda8b42a6a8aed3cb6018636758be3051cee87758ed5998aad924516e34c49319b58cf00000000b7f0c29548e1c1244f0caff38b285b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d6a32076b2f85398959f54218befefc3ffaaa3b7a7272bb85ed06768, 224'h1ba42ebb3927b3a77be0bb8359a91566728fb6b79c206bf0fda960ed},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{278, 1'b1, 512'h1c0e382d29f7ce824206c57f19794f9e8abe01e6af45a57dc9c01184c7b956aba27c6536c48c0951e2540bf566ac000000006db962ed4d45bf0d0c1c6c806b4c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008707126e07ab9635cb48bad9e9b03b432329ee158b173bd8753e3f44, 224'h1214617e1547956f34f9701d4a73958ffe91d9fafeb8b28fa38516d9},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{279, 1'b1, 512'h92cc3187d3326341d51f43165add210d496557c7a27669692c21c2912bc85d13d22a15ce9f2dc8052f89cdb3444fb400000000da250c8d1d81c198686e0c62d4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d22d8e4cd378fced312d893e6b3b4c0904fe2932eb805bc0fa2ebce2, 232'h00f0eaa7c6d10fba23cde05be6dfd7a12ca7782cbe2639f12154009494},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{280, 1'b1, 512'h0ec91d81506646053327c352b11803f36a38ba32d940cdec35246744477eb4c423fd81dfe4e728bea623290a65646d9200000000f68a3961185e3a1eb3a74496, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f6e406ee55ffc2a61f2adb63e3cb19284b1c067c128cf445b68dc259, 232'h00e17e2c98588ce6cab01ac7bba1e3ebe1b45266563d1482c920ec8e8d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{281, 1'b1, 512'h290ba1c9dd4ce7537613a8092317a721e35cf33f17d8c82bc20a765683871857d7a7f0f72e659928158b11760b339f16fa0000000065c91469026a04f6e368f6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d91613f7e2f1456d833f2c9aac0796366079e92f2e30985440a29409, 232'h00e67217bd2b578172b9f225c7014d6cdcf875cde0428e51551b2959de},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{282, 1'b1, 512'he9caa5454fd145db00275838ae34244a94ee61a025a174247c1b8056e6959c7f851f3038bc773457c88404c0dd497580644500000000719f683608f5718616e5, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009d0d161352c289f9b1021b88c467cdd1e6d384e3e4019da7c56c492d, 224'h1c4c4be4f3c9483b5027b5fc7d4729cd74c3b9cef751ef62d2250199},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{283, 1'b1, 512'h1827524c50d2a178cca81cdd33a0be182f764450e04af569ce80811e55ddf11bf9b04675631ccc24d816b26e407df93f288bae0000000040fb10fffd72f8f6b7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ac98a4d298b096e78461602120d1660311fb8ab1f18b46eab3da4d8d, 224'h56ff93d698fda5d8d01a5916ea6d348510f2080c8d784e801a83be98},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{284, 1'b1, 512'ha5186acc06258c75ebd6c4985b00ae514a23405ece5e1c0a51122b5727c5b17a8adfca46c2479895b4121c304b5b2785c72c06a000000000ded1a008316d23dd, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f61ab89eac55f6224381071c2343df902170b58389edcf7e5499cec4, 232'h00efdc8158e8392dfea1c55c5d62ae7b695f822a6407ce52c3dcd2f823},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{285, 1'b1, 512'haec77ef7d501e59ceb458f4b03194d730583d8282b6bb01ce0b0417143ca15c2059e8290afa26d6c1e38502d0b895bb4cb182dd4cb0000000097ca7caccc470f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e73556f65fe40b2599b36abd679dad75fe951f32b7771ee6269b7470, 224'h687fb6342c4bd2f3a215c0405941be22602297164fa9115fa97f58c5},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{286, 1'b1, 512'hfac59bb2cb17756c53956cbb809fb1dcf8f30340a8b21f7a25a1e6b500284c29820250c5c8492ecb2f1c5906b55dfabfb8c47b418d50000000000efa79a0e20a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b1201494285b63e42b59ca8bd67bb655f41d020487c6d4b45c5268a, 232'h009528c4ecfb75628ecbde99aa0a130463a1df91b0205de0b726fe6fdf},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{287, 1'b1, 512'he1942b44674c9c247d1f5857111e24baa87afe02ae74ac9d1ac122c10ced967b6243fd3055a4de1d50b98e24831c9f613d767a3060f7f600000000e5461279bb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4e029b6b69d41ffac3c9d46c79604466fa42a7a66a6cc873dea2f554, 232'h00d554c422d03c2642848e99400aaf411d6ec81fa0eb9b43c4c0bceb1b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{288, 1'b1, 512'h9ea149f211e7bd1f624b20fd50fd2c474d627b16250fb6281c6bf57af0b868f48101c656162b5e1415c87cbb7a685fd752937f97cf58a424000000009deec0f0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7b98c9dee7ac12a6c2f59b20548a86cafd7775a15fe290d48484dd44, 232'h00e6690c32b6b1aec825cff9d2d47a1bf5d6d20000983397bf48c04ce2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{289, 1'b1, 512'he2d392cec1344167d947974fed90e637c5f80aba4fb00ba57dedea9f7ffd1b0404437d90e50f742cad5ed8b82bd136d13319934da1f04f50950000000059c93d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed3385dfe122f21259b55028c6ba2f9ac94594bcb5847b764677dc7, 232'h00b5a12a3f4b088561e1a007e4f052bcffaad05b5e727f3e9385154063},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{290, 1'b1, 512'h40195fbc1bc4b600980e2c2b763857780d875bf68fa15558b038d9333a6c76f3aa4687e0325e29c3945bb8ac11ce675dff92bd5dcf0efe1264e900000000cdc7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a3fe5bf1eae043dec8021e5bc9090fe8d5911c1d6d5a5b98b0f888ea, 224'h7ed55be1e9ae728fe954d34c3effeae42d5f03092d7eeb0710bf1d5a},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{291, 1'b1, 512'hafc1cfa16e5549a03769a98e0a323b3ce3d8e3f316cd9f1007e4366b81a3affe3acb663d6a5d6a6857c736ce28eb85c432aad5ea98a80abb0b973c00000000b6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3e6573e0dc060ec88be161ecfb2200c6f7ff5127a13820bbc4602a54, 232'h00c852d88755d4bd244f0acafd418e499245f2e6417dc8be725143b1c9},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{292, 1'b1, 512'he47ec71fc0cae21e08260f64fa9dc1a4c99ce92048144beeaf932a124c0f87a8b0db214e5424891f30a4cc0311efbb2d49807cc31733db9bd80f912800000000, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ccddf99cfb3ae06c478e62b499cdb2e5a98c665d5fd323cd6733f262, 232'h00eb3b93b35ddd9262e3174aaa32bcf46aef4becd9916166fa3d7cb0b4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{293, 1'b1, 512'hffffffff149aabbf287a78cde6477453f7f9c2310cd2d58ece43bb07019c69c965ca25e8df7696c97ee4ecd4966f7577eb41a60745d031a94f5856e1a5f95aa5, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h088d461e34993c86d1520bfb3a90f1190e08868988bc623cde1eb879, 232'h00a118136bc47181a4edf9e05d3db4eb5ac73da50a95b751e48939be39},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{294, 1'b1, 512'hd5ffffffffa5bd8691d54adc06abeae7d4857cd52aa3ebae84fb391361d804a381d15d6fabbedebceef14c94b5bbcf1560bc8b97cd4c4accead9b453f6d27746, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b51bf389a898407322d5fe142ab2f81439005ab9b4ac3f4031c06d43, 224'h5930035a00f6a1bb805d8c7acdf42b18b020a9426ab7e2ce41f3694a},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{295, 1'b1, 512'h9481ffffffff6e35dfab283e61e8f9a49de1cda44cdf1e2680292ded627b16d9b566ac057cef4c3380ee126c020a6ae86ded132faef613440c54185ed5986dcd, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h565c6827c8f18daa21a6b1edb8af81193e8e391f3e8360b346c7b98a, 224'h468b8b2e16c51e41e26651493e02f0db3af5c9981edfff2991d10599},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{296, 1'b1, 512'h2d8fbaffffffffb42e8498ddf2697ff4a2223fac0c486f05f57374d84dab9e8d13f52f6c898c8a7a74f2d48bee3cc16265e12a6dca3bee77c0ff0ee5e9af7e49, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6030ec07ae1cd991dfbc6b48da43c6240b5bb8f7fe19832df596754d, 224'h54b93d4ae52e4cb7eb969a1eb62f0be395d30a43e7d5736df6b508fc},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{297, 1'b1, 512'hae17b907ffffffff72c833830a0827c91ae711b1704754016d3b0ef4c8367a7e93d4ba6f63e6bb8d572c24bfdc55da0d39f5fc8def9b04723ae25c1b82a3ed86, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h75c39954f9f95618cb890b1a90b9e4fb5b8cec968f8968f53819d497, 232'h00cd93fb7f8aad56fce1734c81229c6b1845635631209fe4d35a4be97e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{298, 1'b1, 512'ha55ecf9029ffffffff0b0266df6f2fc70941d6389583046c5649a1740aae64600c31269408a3fe8dc0975b57d60cc95053b7d311b677bda6e8a0d6792e328bb8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1fa389d2f4e586d5c1e9fcf34b56ed6d35558714d565a61924c59edf, 232'h00ee1a1f53d0f65e00c6fccdeef35566e3d3cbb5b910127d0a40025318},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{299, 1'b1, 512'h37837a8407b6fffffffffac5686980dc2ad1a556be4d1fcf5dc000a18139c2322fb6d35995be1b96f942fa8bcb31b6d4c0efcdb2febaad183b00f4967c63c04c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f1ab78cbc3c60bf97e583ab50abe7c96996b2af0c71e1371a94f9235, 224'h21ec7108be398f859f8f75a8b9b527914685c5f3c1eb26f9b0d44414},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{300, 1'b1, 512'h148ae8a9d1f212ffffffff9007e49461386bac4123a9f847a6901d8d1508c822348ae29c100f38e169470e9a05b8cd6c780a06d49e062785dbdf1fd4cb89afbb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h50e0e423fca4194680ffad95d1e5df534793d5524099addfdaeac0f4, 232'h0091c4495ad79929332b1ca31a3b7d4b94a05b544d029f8df64e54d170},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{301, 1'b1, 512'hc17991fc38743c0bffffffff12be8c0818873e8d65ea350547aa4cdc067cd0a4c21e1d9387ca3c60306f95160cc1f85a08ebdd4f3107b359483b719f5b9a18ab, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5dd7d39e95169cefd77a5a5dfd435e2a879576faf3a845d266d402ca, 224'h63225084b9219b15884e0cd665aca92ef1f4b541987b98cbd03edbfb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{302, 1'b1, 512'h45477dd24fb261b2dcffffffff376705fc972d1fc0eebc57960e96dbf0315340601ad9582193434f8cf1ff955cfa9a803a99d9465ab1d11337155273e65b2735, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00902fbc7eed7ca442c94240c75323db9f690a84817f824bbe12c2f9e9, 224'h12e49c4ed88909344b61c4eefeae4aae0494044bd01653e66dbc480e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{303, 1'b1, 512'he4d30dcc9e0b433fac32ffffffff83bb0169390c4443bfa7b7bc8a7c4421fb94a64d266b35ee622ee92a194a9c369a1bdd0961e4047a4fc3ed632b51f01547c1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h16881c4ae60f32a6b81d445f7bb921ce4f4dcd349695efe0fc94d213, 224'h06066332f61edc98a88a21a42f26e912c99c5471093aca9b1c11d54e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{304, 1'b1, 512'h8f46b06e493783b6d3209bffffffff5f263101ceb63bd0313945c63e59a123011230ea2a874c147574859882f49e6fdc842cbd97843daff440629f6a58573ee8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3d0af397602fc0d18d8a733377cc3e596c143f75d6a9d2c62c99f327, 224'h30ad8bf0bef3b8a2bb4158db621de4570d75c5fec7bb8c3e78af8445},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{305, 1'b1, 512'h34de554e38945bbfefa7cde3ffffffff7b63c616e7853caa71db174d8c61626ec0c2d1fc20cbd176f51bd580fb3d6dbee8b1319ce824b44fd820e94589a562ad, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f95c0fbf6c90b300d80765d7a5902ef690d4dc9ae9acd20a3a7b6d78, 224'h73f3ad08dadaf5c5854d351d47e4ec328013eb7ae9c7e83e110024ad},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{306, 1'b1, 512'hc80ad608a993f311fc5d85b14cffffffff76d81aa75f097430416ac8d6d4e8f80858d995030cfd10467787a708fb59252ba27fd5cb768e2b3cf03a351aec1402, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b324aec4420d11a7da67d287198abbaf2c9e6606a231afa0924d5902, 232'h00db1ed6b990f65ebcdb8c5bc38c7e1b83cfc8f8d00ba4ced39bb565c8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{307, 1'b1, 512'he9f4410a9857187394e0dbde1bc5ffffffff22ae4f317b16e8c82ca5e8ed1488b15705fcee61951d122b9603a8b3744eb429a850db99537b15bdee559ceb17b4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7c2088076ab28c40279abea3fda0a2286e0afe963bacb5f70ded6555, 232'h00da358407c1cc5c2e776854500f44a904b2624ab94ce101fb2b326eb0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{308, 1'b1, 512'hdbab4c37e253fc1deaa9e71c035737ffffffff6e927ee1da438de0d1d5152cd6d0549d2b8172bfeb94749da7ff020aa760407bc5e12a5a099a45a301588b62c4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00abbf69e074a39e167d6c4a61fe0eb2f42a42afdbd840f63ddb3e057d, 232'h00b17ec9b01070d7d8825969bf5f72aa047fb4557bf4525b683a2dd061},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{309, 1'b1, 512'h2ad0f69e7f2e5efe8116b4b576a322e8ffffffffd986d354530161e2776001b50987f4eaccd1eaabb1c1d4d6c94e4f7460ebae1ff8cbf4a1df1cbf4a3e01348b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h787af603539b58520ab74999fa2fc8fe90ea10f3c1b16a181fdc0954, 232'h00fe25a9b16e66aa1c50a59042c1ff0a85e2f4811a8d7540f83a632684},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{310, 1'b1, 512'h69e08e9fa0546aec130be51f245d0daeddffffffffd8d24508cbc6106330bb7e4453fa88ddeeb7a8b80db338a7f66e078ffe0ee91d6b432c2d52b5a0a15f847a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c6fe299f384a978be18fd5dd2e94ca1df248cf17819c95d1b317b257, 232'h009c2bd111dd41fb56a9ded5ce44cf616c3e735e868a1b19d2575fe8ec},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{311, 1'b1, 512'h21e7350eaa2b2a36fa211d7c6b144fc87b5cffffffff9c3a4d277dd4c34a428a3b35dc4d8c1840740df3876a387e6ae3c97b0a40325ae41007bb1de4338ded6d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a68d4678ce9e0cee7ddb75bf4b5fd162ced09c1bdc366336181e4dcd, 224'h2898aecfbdfb33e6be1ef59a20f307729c9954ebff5f119adabb642b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{312, 1'b1, 512'hffde6b2d174d86702f3a46946c7167cabd18feffffffff2df58cb555aad0b0df043b0c01b91bf2ee4827aac1d987f3174e1fce7921c831a0b0aeab1ad1156fed, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h32c28f726d79d4610f6382c329a3a955059f5876ef343585098f40db, 224'h20d7df0ae11f3909ffdc54b12d05bd294505ab76058c79c61dfceedd},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{313, 1'b1, 512'h55260440dd65e8c48db54c801af143d639f08a95ffffffff9f03419e88a5145c37a3193cc07c160404a9b7d489aa324965d89fc40fab65a71fae34c56afa395b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00900b8cb66d0e2bf2f0c4bc3bf269b521801e888ff17c5b8286409ac2, 224'h6a0e9736ee8a570fbf7686630c9dc2613cb084c645100b3924b2b8f3},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{314, 1'b1, 512'h16438d031fffee5b56365cb1a8f4bc19eb046a111dffffffffc16998d3235c27ddbfe7f1e45105d70ecb963cf511b0e09daa505bc426260466ec6528fd48b88f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fad47b9ca7acb94da34cc59586a9a42b95a52d809e3d5816cd1f2af8, 224'h42c895f05a25a443ca32a070aff72225114b557734b966293b657eac},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{315, 1'b1, 512'hc0635b12b9164d0a9480ba133839afb60f79f6e7fa22fffffffff18d9363b5c503a5ae2f4cea06d8c5333965149a2cd0ed0491d1f9c8cfbf12fce9914dc22f30, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h431e666843a0d5e131567ab13ec0accd1fef8d441e96c4b8834d4e40, 224'h0e7a8bb3cef5a676cf4148da42b61457cf9fd43c8a33241d4bb87181},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{316, 1'b1, 512'had86d31823a92384efee57d7fc747fc6347312c57d7e61ffffffffbad8263d3a80dcea096adc61333c39ceb1a06bc016fba8beaac8adc0692127ebdaf8bb65df, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h41327e3497a615192c697ae6a6f8622ba493987f617613e76d134f26, 232'h00e2539f0d6121b27d4f7177714ea5ead4f4d49284243e3ebe964f9c47},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{317, 1'b1, 512'h155ee257be62746434e431f20477a5a614b621ca050d7f78ffffffff517e6eeec93db0df6b6358b1f45efcb67e7b201fe4b0f7ef4fe49aed869621bb74d2604a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h37506ccd77f8097e83d63c3d52af634cc0fe98535688d962b0bc3689, 232'h00bf89ecc570436c2fb85beef396422626cf03f7c2dc16d46951104496},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{318, 1'b1, 512'hde8b1dea4af73e03d31712528653ece2fa048092693f2106acffffffffc4fbe785cc6cb125a5ca069dadd2dd809bc3c6246bc299c2bd84aaaef1085a561dd79a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c97fbc5027204b811f4c250ccab741e22876d1a8f8c6237ea915ca38, 232'h00c51cefcf82a303935b015f0551af07b94bb2203e2bc7cbd34520a35b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{319, 1'b1, 512'h372064a97724ffe3dec873aaa5c4e830fcd9ac84f1c4edb9a372ffffffff621efd798449ba3d7c009467fccb63c6e9a825df2926734122b80e8fc9a6c956351e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0c1f93e9bcb1cbddd0508bda3dad7a96dd09f1321136708b586a1eb9, 232'h00947ef9a508ba969b422c1d8e16a82e8a06a0014afb73bc1f1b6d3a31},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{320, 1'b1, 512'h0a55bcbb94c925c397b334ec37bd5216789d87fc6589738cdccee4ffffffffbca7bb2e94ddb13839ef8da502b39ac80f25abca143e0add021592ea7a36ce83ff, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fb0ca1572c10b3961e9539a9423a55dd08dd991fc04e13207b801a7e, 224'h7c9c049836e1566b889c94416c04a4a861f3573de771be3ecfc0c6ca},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{321, 1'b1, 512'hef503ce85b5b48ef35abff5d47345a71aa715f5e8e1568c9721a78ffffffffffe6124c567f2fb5b5f476271da455e079b655dc8c9506b65d9e3c60892984e8ba, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h762764cf2163759dfcf7863b20849c6deb57808cb208479814a243f8, 224'h7b41a973df219ea717a653bdbe27669bba57fc7c7afc3afe9c87d62f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{322, 1'b1, 512'h5f3afd4f98713d775d93b166838053fa503faf72cf3c00b3c57e0fe3ffffffff7b74af7667db987c9c205466e00679714af8467254f2e441ccbf1bdb9daad40a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5cc108138881be0cf7035dcad94db36063eaf148d24fedfe44723e5d, 232'h00d11637a4eb1e2e438593eda38970537a05590b3a9a5054d3afc9e9bc},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{323, 1'b1, 512'h9e670958749c5bbc0cacb1ee6c38e71eede821d75d84cc2fe1335af9f6ffffffff4e9613cec31f535c4c7bdab269d70a8d4b3bdffa3065d91435a4237cae96da, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h531c06348905bbf16d85b8eba22f5d5ca33e490107ea979f6f322a65, 224'h0109215bf6d2afbedf4efe481f704963355f09f59e1977be330972a7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{324, 1'b1, 512'h1e77a725c36046bc3bd6ca38747586093510952c0a3390d86b508479c0d6ffffffff25680ce9cd685ebae3cafde6315263f7cf4ea6117ccf870d42189ba3abb8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdc683a5e7cbe5df332c85af8c33d7ede2e272dce6b40d360d666acf, 232'h00a779a6f1fe92ba3f799595289d7f37d47a1187285d7636330a217a7a},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{325, 1'b1, 512'h59f9626626a34d5491d567d0315894fb702c1d7a2ec677a2b595a772b20d8effffffff20557e965f33f606242a59aea4cd565aecb931664e51fee93a92ccaab6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70ba414a666f89e84064b2f9b08d500c6bb12d0a5ef9b23f4fa46ccf, 224'h43d88b7e943fe8792ff62ed462ea308d28f7f03e4dc59d6214f30507},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 512'h001db8dc4aade36062b6ddb62bd342923f537cd35c957b47803909be234a3b58ffffffff0b537f24fbdbfbefce08b061b467fe60e7f86531ed3f54c6e29889dc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h126507852f3606bae527749982c5b303870cbf999d2f0191f5fb7c62, 232'h00f4c92989775dd4183c62fba423e628fc124db1718647a69316e0614e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{327, 1'b1, 512'ha05bf269c6959e1000f754963c2ee746346fac0d57bb119d3cecfa3dfe702fef2cffffffffddcffafb72da48023b4eae3593eb7c3c2d758c1c6c5e4dc57d53bc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009342dbbf6c92387699c84cc0f8b011690c072f8f067cfd5de213ecff, 224'h09326ae7030d262085de892da4cfdbf787cffeaaa71dfe0059e28b6f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{328, 1'b1, 512'h9695a59c40d735b329f1f9c2ffd974ea8e66af6c65a1f7242e1eb02ea6721f9460ffffffffff9327209276e0633e07c96c9a2950a09411d1eabeda48ba90c8c3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1e6e376f2143d020848ef2653aedf7123e27fa8c67585655e7f9e5c6, 232'h0094c8ea3567ed7726d5a145f417ba44bf7afd586e38c83748dc227830},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{329, 1'b1, 512'h521abe64cfe7fa37251542760a99aba478c8b79a5eea4ba1fa859e6dd8bf23196e36ffffffff157c00247c6e0a683044034774f96f67cdea42afc9ebe8d78be0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0099f67a076a74ef92d33cb89e39944423d6b60d6479f22a63c2b2e6a1, 224'h1cbcf7baa7702cdc175d4dcc3d6a016e90046ebf74de51bddf41deac},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{330, 1'b1, 512'h56f7dac71cfda3cdc27537a7fef1026211918d8041d79637eee4bf44f6fda371a67755ffffffff1dbdc9ce7d24880544364cd8cd5925c287a256383c78631a0c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h61ec8a8a6ea82e842202f327ca3e5971521be13c6dc605e779fa9b47, 232'h009f87294c702676ccab8a6b31aef5aa104139da7cbc69b1a6d4d77a6d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{331, 1'b1, 512'hba44f1aa7dbd00300b9d114936943eb2585a2ca6cd8f11fd68794b5adabdcfec1919ade7ffffffff099e11a571237729c09fc81d86398317874c3722999b1875, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h467ffbd3372c95547537212af707e412919eb3731ba661a2f20eca59, 232'h00beeef3b4b325d5004f0dbd99a735778db53e0aa381a069fa68f00852},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{332, 1'b1, 512'h125406f9b34e4f63c0a2288bf6166292074a0fed2b2c47822bb885520f2db3e2c58186b926ffffffffee3b259d2c85d9ab10b9f10f7f3cab27a8f528b4a82ad8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d4bbeb81922f0e5f10d637a48dbe3d80cb53524876821dc2fabb3457, 224'h23f8ff0919d566e05a26ac97d51bdc79ba9c920e2d6c777b8d7cd4e4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{333, 1'b1, 512'h46943ed052f77d2e9549dfb8b9a4c779959f7b0a78d6bf2dbde3be53634e232d52a793b7778affffffff162f29721e93b2c9de6629fffbe68596e94b26703923, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c151ab28d7a23986021cad0f2f937b61c4adab21acf5081cade56585, 224'h386aa40927cbc45216568b23f6a4c49aeab525e94b074b8ef16aad64},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{334, 1'b1, 512'h2b88c2f7b3ffbf92cf6698268ef14cba56c268701a73b30436de1465b85a572363de2fbe10e2beffffffff9b6ad94f832c537e1e40dfd29f836574fecb7dd074, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h40a4b6106960c1b249c116d539c9ab27f992f0c1e92d8e04a919a749, 232'h00811d34da166b2447a2da0e3821cff12cd47ae0fb273fb18df830d179},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{335, 1'b1, 512'h4e29d13bd24e9f13d5e31ac769469a23d44278a67b110f7bab6095667a3a5180bc8124849e31af47ffffffff94e438c9abcb1301833210026c068417d2da4b20, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6808f8c1cf3a051724d074ebdc85fcdc14987324605a81db7591baa6, 224'h026f5efef2c657bc048c88a165f885628efcad293d80a5cf72855491},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{336, 1'b1, 512'h5199a888f66bdde1285c6e1d75e11ca4a6fa67ceafbf32d81894eb60ba36c4786868dcb1384710d5d2ffffffff3d60d7798468aacd9f552c97fa4600343889c9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00af7177ec82b907cafe3ac3bfb0ae2f2a2a8355380ce8b31217fdb3f0, 224'h05282a1dc81cb458f1c556877dc23301cd8f69a5269df683ba1d959b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{337, 1'b1, 512'h7692bad59be557b4e1db6cf148e5f0ff3c273d29d9017b90c8c26236cf78465b335a40716400ae0aaa34ffffffffd68ebefa85c403e0a25dbfeda3354bcc2a84, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4cb87503bde0aca323f93b04e1735f84bc0e101ba8b71332fb40ce4c, 224'h0bbc59dac149a5644771119b00d1d72905e4b080f9aff5d6a42e1565},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{338, 1'b1, 512'hadf9dc5a02f2bf38df234e566f0b5ae3c8b5a20cecc2f8565bb8f756ba59b295004e2ed1807a1e579596ffffffffffac7657366f92a09ca3685510feb2182e3e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ae09718e0e6e7fb0237056f531221c0c93306b426a985ac51a70a831, 232'h00b50599a416553c34102a917990c70c3f9f6ed01719fa9e009c14a230},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{339, 1'b1, 512'hf9db531c8bd06c7272a9ae2de6b4cac8e0281438eac5689c7f763241db7b88b4a6c71d53a3d03222f6195dffffffff0b690ef5a310f733b13a1bda4fe964a38e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7bd61f75610ead312a227d5368e093606a4630663825490b392a5a65, 232'h0086552bb6f4f3564349fc3fb47073c3c28d10d9daf5b9166a82f8a6bb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{340, 1'b1, 512'h273f59b9ed631e0fc10467687508d817c2229d48e45efa2a6783290c6ab048c048a882eef2730e7456b3d4b6ffffffff0369568d9ede46d524123c6cdf78afb6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a3daf123bc8a3e393e8d669bd76c4486a3e65bd16fc390e09b2308c9, 232'h009c680cdbca9d3aa378cfe60481b2e68d3b3687363e6716542da50a72},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{341, 1'b1, 512'he6ded1492cb08b685e2c14f2f11d4bb2fe1601c47019cdd5bb3a42aadbb88f1335fe76ecf455cde30b30e18d35ffffffff921892b8870a2d1248dcd97ed5449f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b782f0af6552a3f30530942f35160c09ec77d06595aceb9da8d246ac, 232'h00f41b8216ff29fc92655527c6aefac0bab839c18525c03316b46a4edf},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{342, 1'b1, 512'hef9ce8e0e84c667ba940ccb1d3317daddea8b9888a2ef5b718605aeff060c7140522f73cdb7670b0e055a2646509ffffffff81c895857965435d4c4421eaaee8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ee945c87a9d4e74d87471f83e4f791945b7733a1bc75fe6738f23ec, 232'h00ab06858d113616b694d36ffaf1736567d3895e005e80f521310b5ed0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{343, 1'b1, 512'h388b354799942c6595ba49bc6bf8e7ca5c06c6ae8015c0f58e69192d96cc60e30696c1284ba98c1b22c5c7f23bf8e0ffffffff15f579e355c7258262f0fdfdfb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h733752fa2b90121c01878170f2019d9c9a4b1c95e82acab18ae95d71, 224'h358eb5d69942b4b5d0d900bb843d79f90af54663b3a926fabd081d42},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{344, 1'b1, 512'hc6bf307fea8c2799ef482911ac86779072e5757f934a3671ad8c5a9e372bb2ec8d318ee3bd0cc4460f9050c937a3409cffffffff81c81c22e9468fd07ec09f55, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h72fa0cb38863c06e535402e010bac709ef4beb0b38118c7b13308e83, 224'h33eb21f6c081afa7db62c2f8cf78ed1982cb762a130509bdb53f1774},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{345, 1'b1, 512'hf5f21b002be6b7b3a605b3bcc5a3a12aa0b905565d958028fb8c44d8e5182b6ea4beafe63cbdd96daef63b98ae46ff91bfffffffff3ffcdb29cde67329851fd7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009277ca6db735f44bff16c7ce43ad45707bc6a6b451e64532b86b54af, 224'h433c69a072349f3814c6366418d3eb7fb05509ad099afeef411c6e11},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{346, 1'b1, 512'hd88d68932ee321d611334d87de84ef4240025f9d0c8f11bd9aaea2e7729ad87ab0ee66d229b2eb78221050b375a54bd698a2ffffffff0967dbcb983a8f09417c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h37e05ebb376ede0d3fc7528f19dbe4a38e4f310295058e2173f88900, 224'h4f8d5ca627d43c54db6674e1462d12c42603cddc6f3067307ab04d4f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{347, 1'b1, 512'h611df311628ef69305da2acf952b7289eaabbf389dae756f08c459819db39b7133f02dd126e0442f19bce8ee83cbaabdcd974cffffffffb7195ff14e2d445864, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a419d09f64d28e4ca617187790d046e3b29b87dcd6007eaeef08aef0, 224'h397fae569961478fd7d075a30398a646d95c00f8171600e1ca2335c1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{348, 1'b1, 512'h4f34828f9520f17da9e588884a26df5ab85e8456184bb19001abc926a180c32a112ba4164e81d69b8fdaaf3c60619a7d1a5840b6ffffffff8748db5ab09c4a64, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h05ea0f04e9b4eb3b62fcf8f1f1d120e58a932ca9a04e8c64bbee537e, 224'h166633a3c8d2b5c6246da69e069f2f09a7912efc355c405302b2984b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{349, 1'b1, 512'h4a3d25b54b17b001046f323462e30475caa0fe686e8fa4eaa3b0cbf604de9812e2cb4eafbbe44222356c1e1702c09078e7df08dc98ffffffffff06067e01ce41, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fa2a6265e9fbd317fcda0adeac307fe2f0a94afd6303c91985d84d10, 232'h00db93f0201284b5b66a15ea177f34c27c6d80479c18db44f386e85d37},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{350, 1'b1, 512'h6a763ddd1f348cae57162f918abd67d536a03431ed29721e179403366c3fe64f1083d4a64cb7a9fddc7c5a3487675be4078be3b484ffffffff2d5a70dd12c49f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2d58c2d0cbbe7215424b943006dd56d23159ea10140569dc22663bfc, 232'h008d9bdec0639a236e95fdb35dc2ce3d63f7d5447b6dd3d95227fba0a1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{351, 1'b1, 512'h0844602883dbcf60972c8b943b5ea020ccb0d19c82eb86cb18d4225a79f97279539214d6e3df6ba6af165c9cd95b8b67a36b39bbd101ffffffff5a9aa9794dd2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1bc64aaf83515275fd3187a18d3651c75ce85b53f5579ecf5f190334, 224'h2ed9fc723bd723cd4c8b62b7968e5f058d25aa6f6bb45e6b09337793},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{352, 1'b1, 512'h73672c1037e14e2ed10a0928e8938944667e83879d16f2688f2fe0087494b9f496471dd4e27f5cfddfc4b5efc4e7fcd511d2f67ea879f2ffffffffaebc4501e4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h240d8b05889274d716f57588536320775afed824d79f41f32c35e728, 224'h25031a073d638165f8c0b46a28e008f1de9fa0cf726d316269f669d6},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{353, 1'b1, 512'h1c28cbb7dcfe2b79763ccf8ebcb7939ea373f7751d8b3965fdcd8b62e8360f619321855d0fe872fcbb3509f48c195d96b1d765983c695686ffffffff51d7cbd7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fb2f81bd4e22230c0c95a7a08eaf9a668f6b5c6d32bffaf538bed19d, 232'h008ae8c126b3168129a720a674fa4dbb81d94f4a3e862b834ea328ed4a},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{354, 1'b1, 512'h823e30e3f8bce86e5790d073d931eed5a7ab1f52fdaa4a2522831c73dff05fdcc91829a51c8c0c97c24def713b52643ab17a700ddfa0988740ffffffffca2992, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fdcdf3940d5b9b3841fa0ee667d4ed9ac74e0cdcde9641270f2e658d, 224'h3167f2b6601b737bc4a700dd0940ef86107eb57c39efaf6b3d71fd38},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{355, 1'b1, 512'hf2104bf641a8b485448e73c4b7de7fc4ec1d3e06eae0f264dbdadb0d514a7aa2ff1567a80e8156c2bd97579eb1467c0efacf0fdd1166e87838a2ffffffffc8e9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h46408d1ac74a5bd03c3fc08685f2743eb3f7c42203f63606775a4250, 232'h009813e4704b565f94e563a653a9d4e0310ebc7055729f89ca4b02d9f0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{356, 1'b1, 512'h3db47a2cad8a1c43f31ee677cef231cda0f3853901676c1732771602ccdcc294a38fb8df77d5e6e5737d4c8e05953aeb81edb39a25931717b3c154ffffffff9d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c9096071c92973198efac69d6b3912e4e14248bb077602870c543cf2, 224'h631c995cab8f0ccf5e3dcb30d4b995dc96d2573facc6ed9561cb9d93},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{357, 1'b1, 512'h6becb022ae22ffc4efd852cec1259abcbd9936403db48920bab66dff9bd34bd1ba5c30d1e8752af80d13d9304dfb864e834181cff7e8be9467cc3617ffffffff, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b55bb2da01e99b08f64dcec6d6d746b5626aec6eae2378fd1db72107, 224'h07f36d4edf6c8112e2a6b9665b19605f41c9449a7eab7839d638ce10},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{358, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e630949b06fde06a763cd457fc1776a006932c0fe08131f44aa1ca41, 224'h3de7e43d3671fa00db71d03e7f4d9f80b0d6d7edb695032e09b93d44},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{359, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h078e4d1a56e6f485c785d01a8cb9bb2ef5c7646fb1e88228abcf5e01, 232'h00ca1fb26c9366cd918628033dad9518a8f8a9ff4a513c6605f5cdaae9, 120'h00e95c1f470fc1ec22d6baa3a3d5c1, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=120b(15B), s=232b(29B)
  '{360, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h078e4d1a56e6f485c785d01a8cb9bb2ef5c7646fb1e88228abcf5e01, 232'h00ca1fb26c9366cd918628033dad9518a8f8a9ff4a513c6605f5cdaae9, 232'h00fffffffffffffffffffffffffffffffefffffffffffffffffffffffe, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{361, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h225298c3aab4ee639834fe16c42896f6478f3517589064717d40959e, 224'h72881bddefd6ef724fec33f92c92d4fa2fffe77ce20a327845b1201f, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3b},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{362, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h448bad17b638f55372b256c6717ac0fe443c20af133348be8f728577, 224'h421c701ae6015da98a2ec4140122091588c013a74fd78b3814c981b2, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{363, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h146e29fe57ebbfb91f2562de124e62408e6c3e951c96fabb83d243ca, 232'h00801067848d29410a1611656866e3cececfc569091375b674d7e4d167, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 232'h00bf19ab4d3ebf5a1a49d765909308daa88c2b7be3969db552ea30562b},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{364, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00fad98df6a5fbd9f3c023f2ab809c57c72de3396d1cae4bc35d78d8d1, 232'h00889e372a90189ece8fbc690fe3cdeeef38ab12ffda721f32f849ae50, 8'h03, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{365, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00d2eaeb6be6b5dced48d595b95f73b069f49a078572c74dbc557fa25a, 232'h00a6388c4362e6aa12ab9c1350cd6789d0955445d9198ecc3a4618da73, 8'h03, 8'h03},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{366, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h2df6ce6019d77e3c6e04908a3fde5b8833f9c493bf3cc6568e3d40cb, 224'h0ced2e9cad2ed363fd20aeb9983bcb22091fcb559c1f6fd538a0ae04, 8'h03, 8'h04},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{367, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h2df6ce6019d77e3c6e04908a3fde5b8833f9c493bf3cc6568e3d40cb, 224'h0ced2e9cad2ed363fd20aeb9983bcb22091fcb559c1f6fd538a0ae04, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a40, 8'h04},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{368, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h0093aa938387897826db23b19903c58a32f8269d93a5366a7a673e30da, 224'h27ac5a515b7081cd74bf69528114241728da26ae6895e83fea25bec4, 8'h03, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c6f00c4},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{369, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h09cdd0119a392a271c4055fac2fa71fcc678b9c318bfb90dd1ad0ad6, 224'h4dbd418726f0d3f0bf0cee7a1b366d9711793c839206e6205c416ebd, 16'h0100, 232'h00c993264c993264c993264c99326411d2e55b3214a8d67528812a55ab},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{370, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h008f711e9fbea41bd25aadf584999926a29c2801e7dbb2eb1dbe0d1586, 232'h00841a143bdeeac9969be87f57b4d71a466b2b6aed24e854b07570e629, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=56b(7B), s=224b(28B)
  '{371, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00c288ddd81714a9e766b35a03c835fbe1a52c540b747b11ba3ebabdcc, 232'h00b26bd049bd3088b553162261eb93ab5a75d873bfca8122a229e2cfc7, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{372, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00fd931e8f08b12ca82a6b050e2c281b0069258ac851131008f9c2853c, 232'h008beabb4bfeff98be4ee23f90b552ccc38a72976bc71e7637dad27fba, 16'h0100, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=16b(2B), s=232b(29B)
  '{373, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h1dfdd350e45903ef44a28acf73999a22a706a589a3dd20c051dbe4e5, 224'h41c1021ff3e9646ead3e9858c9c1bdae1e1532b69b2ec52f8546f573, 104'h062522bbd3ecbe7c39e93e7c24, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=104b(13B), s=232b(29B)
  '{374, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00fc06e8424839eb95203195f9ee12687c790bbcc9a740d40c1bbbcf66, 224'h0d1afa473637d708952954a18067b4cbffe584e9e891403541c21fa7, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c29bd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{375, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00c847d6757702db5d47caf6129e865aa22d6b55c545f70ce7e7ad0eca, 232'h00f69bf4c624111ef1ce92e9e10d126f0ceda9851dcc53993930324d3e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{376, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00c847d6757702db5d47caf6129e865aa22d6b55c545f70ce7e7ad0eca, 232'h00f69bf4c624111ef1ce92e9e10d126f0ceda9851dcc53993930324d3e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{377, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h61c0d09fc40dd59a7b5281af54fd4db8819997cf31212a4b35cf6078, 232'h00a55ef14cafacd57ca50195aa1962aa7d01f7595d76d342d83fed44ec, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{378, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h66539275c7d5ae5dad2507a7169c48a9cff067c4d6afeb22561239b6, 224'h12eec9a7e63d602cf87f3581bdeb19ce994c48b41079ef8186339dfd, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{379, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h43a45adf3cd2a866e01ec45269f604af026a4483973cc4356b473966, 224'h2a8403f5f14fcd737d2aedec136a534417e0d19e1b98d53944100d0f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{380, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h2e55f92435ee396708e4805e3a2c4c6152c69e1671e9d6387c56f58d, 224'h3b4a173ad9f475448586ae0f531ee07f15553eba9828b2bc8d72c5f1, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd543},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{381, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h5bc1eb0ab6349146bf13d2aafd9d44c909397d39c12371ff7e56b126, 224'h4c7f85004a22aa08c93b7b14c06970fa19625e671c1fb5b16e8a0bd5, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00cbd2518ae59c5c357e7630cbd4c3e1b836938a5b4bfac8239a9c54fa},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{382, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h144765b9d78724babc4358b229df98e9d64da22724381ebfe41d7e72, 232'h0086e958c2f6779b8ea76433cd4dce0ae4cd300875ac1c7ad218e57a55, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{383, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00e3fc6fee216eb1fa8aea73fc2802709b2c5cd29f99ed964bcc0806aa, 224'h2dfc634b9050acf568963e3996acf0f2c7656a3bc0f091d7aa1adf7a, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaa0f17407b4ad40d3e1b8392e81c29},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{384, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00e57bf59d8236b7b789d45912eebaa69dba563bc790fca99ece5da665, 232'h008bdd80b86d6e9caa2e9086d226614281cc038a2323083a4184057a37, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00bc0f3a2708cbe1438083451163bdcb6579326cca4fdee68ed37d633f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{385, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00d2612ed20fe786484b8955d658200776ec219426479c69194f8c1baf, 232'h00a3af3aa778c1751f4474cc0ff2db2a834c232ec49e9ce142a51170b7, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2d4465a55b282f252f2b47f9f7bfc0ba40ec4dca29f567940b2d90f4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{386, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h4c70cd0aa06d9ee36a16202bcfc891ceb41a26e0bcdde9d93da8001a, 232'h00ab77b507c77931fc7ee290cda7b7af6ad90d0c97b836ae1b65b6eccb, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fe808b87e0e6e76364ce32fde12f692d69dd3b362ef4cf499e03418},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{387, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00efb7722fceaa8cd19162eee8b293b58dcbd0fdd3dcfcd6e6ba37baa5, 224'h659d47ecd7d2b7f65faed3e9a9b554db19e96948a1c5b954351f23a3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00b836c957342d757ecbd2518ae59bb4489ecce8b658ca10e822ecc823},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{388, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h79e577f8303d4ed74c3a19cabe3ec35bd39cb789bc7309335a5710e6, 224'h43cc437d5793931f92eea56039b22088165693a7d9ed0ffc6188aa24, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c957342d757ecbd2518ae59c5c2f4ebdd95caedf61c68b89387f3c9},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{389, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h735e5bc29ee55242a71953f4d31954bc8c173c40bd84017dbc076d4a, 232'h00ce15cfa865a1b3762e61dd24cf61022bb571a5fc8b5d5e7ea80b2405, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d92ae685aeafd97a4a315cb38b85e9d7bb2b95dbec38d171270fe792},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{390, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00ee2558b8b7642287cdeedc8bca740974264a667e5edefe79e7a03900, 224'h5cf362e47faca649cf9b8f6c9214539ef2eee6b86935185c1fdb3492, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h342d757ecbd2518ae59c5c357e76013b79f087e62e58923f7ea5c045},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{391, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00f8b4c378bd5f417b562ae127f39825a2b05770089b7caf9324d7ce1a, 224'h50708175ba245e9c152bff3ca95743e261b6f579328f30680fb6a2a0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h21f862ec7b9a0f5e3fbe5d774e20a59eb3c341b9e1ff215b446f637f},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{392, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h5eb63f0f7b7ec667588670022e2f0b1124b132ebe16c143d6ed24602, 232'h00af2b27b92a449a4edc20267d25d0a238b43aa7289348a1378db079de, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h43f0c5d8f7341ebc7f7cbaee9c414b3d67868373c3fe42b688dec6fe},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{393, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h280ac7f11afa66465c37eba820aa8f393d13c5634022333c7a2524bd, 224'h5c63b1e9ed18115b589b56270c5c3281fa97060f1d30aef465f445e2, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h65e928c572ce2e1abf3b1865ea61f0dc1b49c52da5fd6411cd4e2a7d},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{394, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00cdc63e73d8d6f4f8770a97d93bde4e1974a277adad53d500cb070907, 224'h533c09379488cb344ce01bb29a2f12d6e0b946a279c7f5d47831477c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3ff4045c3f07373b1b267197ef097b496b4ee9d9b177a67a4cf01a0c},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{395, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h5e963ce90708539b001d821b9884f46ee4ba452bfcd539741d8fe838, 224'h4c8dc874329bd0b78fe04e0291f13907ff5723e8d15146c5469d7d9b, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{396, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00aa7f2f92f8ae99c9bdac065e659a4a2a0540f21369383334613b6086, 232'h0094da15e113f211a6e7939caf1f20acc279a3b5b5b0186451ec8603b4, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00855f5b2dc8e46ec428a593f73219cf65dae793e8346e30cc3701309c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{397, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b97529fb4a1e02b5e81d77b0e7909a2fde857a1edc9fa660d600c89a, 232'h00e5a8c9c55885cc20f54f5c8f423f785caf423d77ba0afc31fc16f131, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{398, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00a4b344981d0a826546855d219ab4ab59d3ff330676d93b9553804278, 224'h41370e4dd0de4d096c20881fc35a9a0ff377b5f06deeedc19feb48ae, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0084a6c7513e5f48c07fffffffffff8713f3cba1293e4f3e95597fe6bd},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{399, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00d656048bfd65af83d6dc3f7cb7d240c9e0cdee6e946b15abb13f4b33, 232'h00d61580a159caf9fd87194b7c9d78753e0e00560a208d34c7dd4c6a63, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{400, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00ea6b3100290627d3e5d8a07d7d167022c58e7bdac2701735931899ac, 224'h39bca56a702c508dd51bc96c63967c359e92db790f72631d875e0719, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d8ea27cbe9180fffffffffffffff3a43fa3662a899627950d4eb64bc},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{401, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00912cff3ab4338f1f09b71f909dd68186cfabeb746beae33700dd923f, 232'h00f832461ccff9b83c25754bc1def8f10c5ffbdca0127914cf24184823, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{402, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h6952914ce90a0e65b03fffa7263f04a3f7be03cc6b801e1204dad313, 232'h00f04726e76989b5b0eabf53787d8c9f07549506d128a148a6b4e94610, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00bfffffffffffffffffffffffffff3d87bb44c833bb384d0f224ccdde},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{403, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h0086ec9d3ba7c6d9498069a07761a9d85e04fa21fd599c6a2664e86254, 232'h00c5900aa4b9882b32983c5e029fe6a5578ac818e79acb20beef73e8ee, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{404, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b08c34e9416743b6a3f52c42041a5fc3011f64dffb54875bc690393e, 224'h6a7c67833682e81719f928df55faac24f488028515b26e03c1c9a02c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{405, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h0a07d4a64b42e61096d0b7dd9674800ce46916617159476ecae94058, 224'h6f0b0584dba9d9fb5cda23a2c82e3b28b1c1486150a3419feecc4504, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0096dafb0d7540b93b5790327082635cd8895e1e799d5d19f92b594056},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{406, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00dcb6044f8d2c6e3bab60f13e6da1896e2504d0769c2af824732b5326, 232'h00b80a5437b9d5ebe6d8eb49e70f49220dd3e2c3c7865b87ec98b53466, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 232'h00a724b1fe4251d5b6cfa15eea5c648bfed7732fbbadc9300c8ba40032},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{407, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00dcb6044f8d2c6e3bab60f13e6da1896e2504d0769c2af824732b5326, 224'h47f5abc8462a14192714b618f0b6ddf12c1d3c3879a47813674acb9b, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 232'h00a724b1fe4251d5b6cfa15eea5c648bfed7732fbbadc9300c8ba40032},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{408, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b08c10bbd277ee6ab501aa71141733cb196b74de463ead5ea224022c, 224'h7f68bcdeead7d74cb6186e32219846424a926dec60b2a227411ae805, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{409, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b1babefd03f6f738fc86d32ca245f5db21f67e7bd919079bd735f35b, 232'h00d9ad5e6886dcfc7f2272b98c48a7c43f1c57a024f2f054fc59bb4354, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{410, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h222b7566f26c8776066f2f4065e4e6ac45a306c306aeab8250b652fc, 232'h00bc63004961a554047c03655cea7dac88e573fd45ca4b407b63967290, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{411, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00f9973f688705dc1025beb72663df6f84bda4a14a79e5953d699269ba, 232'h00886f01e609345596494468378d758c618f49e216287d85554af8eb68, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{412, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00c108ca8adeef82f140cf158a70d31f0a5b66d86612b5d4f00e243386, 224'h5cf0f2fa4466eb35279ca99def17864835954a74d12e6c7e8494060b, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{413, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h0ac469e816565a6a74bec821ca20b88a61018a0335199b5d7bd969e9, 224'h463355c73a2d9c51049f7a94509a9ac4ea0165763ba113a30db999e2, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{414, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h662eb328d24fb548f51792b5563ac3cb237f0a65199460eebfcaa5c3, 232'h00e758d13e7b419b417c8c97c4727c39fd373045e18792ad8076b072b4, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{415, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00ae6d9c0656d363b21e562b56f3c85b6d77a6acc664ad5705341ac262, 232'h00dd3a814ff8f9049e4635351d25669b50b51b30e2a5bafc9fce171e90, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{416, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00aa93b40a88f172a1481aad312f4bcc0a7d92103e42feeb986bcdc4a4, 232'h00e62a7c2e4dd34fb7e518630feea54a6581ce5ffaaca7deea3b26d647, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{417, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h42f4cf939e3aa83c2bf17cbe8be930695aed3feea7e64adf6842d71b, 232'h00a17b9dd00589212e33bc190051be877a455622c22adcce8ee098fbee, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{418, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h55a918f3c19077432b22ceee7c2ff87dfe9ba7323c55237ee75f02de, 224'h110e99ed5be3ba0e0306257712168712afaee008163a693b601f5039, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{419, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00bf184f88a452b3bf85edaea150dd770e90f49c871b5020a0a40deadc, 224'h28e7f6a690338ef4fec8847e6f085dc470c64012b7a747624bc9c90a, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{420, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00872f112ce4aa0ff8efe70543dc1c6b0bd14d068bc88eb6436245481b, 232'h00a2aeb521e472e5e1921af16210fa63d3eee42df5d5ff31e6d0761b5e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{421, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd543, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{422, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 232'h00cbd2518ae59c5c357e7630cbd4c3e1b836938a5b4bfac8239a9c54fa, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{423, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd543, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{424, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 232'h00cbd2518ae59c5c357e7630cbd4c3e1b836938a5b4bfac8239a9c54fa, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{425, 1'b1, 512'ha69f73cca23a9ac5c8b567dc185a756e97c982164fe25859e0d1dcc1475c80a615b2123af1f5f94c11e3e9402c3ac558f500199d95b6d3e301758586281dcd26, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h008de3b662a51308a2dc0651a2f50bb3475376e90bb8418256cd791bcb, 224'h0910c5c50a32a24aad84da25559dbf077e5337f3c3f626fb15d376dc},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{426, 1'b1, 512'h86fe1b4ea7ac8e339d04e40087534c61e245dd4a0c22754a0622642bba56de900b2d431e859a36b1a5ff71aee560522eb0d3251e018c2cb6a10b82031cfd37f2, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00dcedb02afdffdd199b47e545e1396a1b170fdf96a10ee4d3add2b496, 224'h4a3c894b80de1bcda509ab58752e0056dc78d6683a85ca9f15c251b9},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{427, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00a7cab432dc7abf269c13632589d9d9cda37482db9e8dcf411c2344a4, 232'h00fb38ff0bea5f81595615608ad33494cceaec48ee6007d4951d2d5bd0},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{428, 1'b1, 512'h7d795fe6a97761d89b35f64e09555951f6ec2a669a9fa03481c100ae158f183e2171e142437d2c3a42352108a22a7e3d797beaf6c3075db419b6f4acca479c83, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h0316a2259370447c1b06f51f6189b033ead956c11ebbc3edbdc2b5e4, 224'h24bda2d065a0475c9fc5ee300f6c4c826b07a740d4990fcc146006aa},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{429, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h00c8a93a8f1b3aaaa9bb8e2d8cc4f5b5033a909b15ad81b2dae14c1620, 232'h00e686820912f295c9c1b31e60c1fa27d8d0f49c017249380f928ecff2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{430, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h3989321934702e535635459d9409606cfc4634c3b282fa86a93c8016, 232'h00c1f6c399ccb2ae5a22e806f1413874fe57cec917b576d3ed887e38dc},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{431, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h008c97232cd430bb32dd89f5155205f6ae03f173f88a1be96a2c33d9e1, 232'h00fb3b4eb539553d6645e434befa760c9fab3d2ae645ced03fe7713aa1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{432, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h72791a86439f76ee409629d923fab73936510ef89349ee4cc304b915, 232'h00ed67c5eedc4a59af13fe80905199de42fbc45eaad6bd44329c7c75cf},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{433, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h24575ff9e5ea779d95644b5ef9affa6727978553df3b51fbc5a27820, 232'h008b2000b4c02a1fcc7880a42c6dbe07e322ebe20940d6ff32a08eadd9},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{434, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00e55819d63e0cdb616676d16d1ad6ca2bb979be94924534dba3fd6f3a, 224'h4dbc47c830fd85e16d013e056b2f0b1646d048cd6fc21757af428f05},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{435, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00d12c22b4ef1ff2de70c6e1a2c18f7dc87dfcfec225cb3f324a76654b, 232'h00b64bd7dd3e3184073acf584bfd33dbc3712a89f201386312f713e1da},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{436, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00c8d06f039201c03995813152a19fe52e3c38cf32b0f13b8d8cec87ba, 224'h449307f7924fa276ac1ca82973d5f55fca7c6690c8581dbbe5500128},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{437, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00a370d277f28e3c86c9367e2c1d7ae07e6b0da333da65ef2780b39e00, 224'h134f5f55e3752543f960e0e7257cffe3ec417b9bc5da3b7557de44ea},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{438, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h2336af69da825fec3510681c716c9b5000b17ef1e6db73707817b145, 232'h009ef59c120ce39e4c83e341af71d4a91a34c4bdd12c92caf4405b794d},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{439, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h3fdb17cc44c9a0e995290a458c2f64b8565541cf56139575212ec168, 224'h5e51c778b560f3c61bc3bf0eb50ff8d34dcb5eb85cc25b4ae6a7443a},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{440, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h1d98253a63b83f0e042ed2c342fd4217c29f990fcd5b5cbb9e51721f, 224'h49fcf5e4d680cdd36405c514414cc47d9731a97c4edcbac7b7b27f89},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{441, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00a0f6aa5f607f34e49af976d8b0fb4f42da17fd1c2b03b8119f7b834b, 232'h00ab5395c0faa4ee5310625d501d6a0af96644040a335ff8f42bad65d3},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{442, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h009a0f67792672dcba4b19899ba2e35ac0b54ca00ca4957270e7a43f8c, 232'h00a702887888511dd12e950eddd239b4a3c423da673bba882082954a0a},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{443, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h4d96e743ac0dbbf2413725a193c7e70947b59501601e337665023ee2, 224'h764ef71a184f0244c0e1de1b729b8421be53bd0ded2015dc3d1f1a13},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{444, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h060ac961eff4e5053f7045b9ea1db338dd4b3a6cce331386d3988655, 224'h0cfc61a43a67d0660fc386efc1b603b28f651885bff519c632e11a8c},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{445, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h3415d0790d9b9ba8ffa82f447a4fed58cce3ebbaf43b68c162495c85, 224'h1e0e20ac93d19dbd9ddd632e5c0910560e941acf2ba5d7f3f2abe27f},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{446, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h2066593be10db4111e032cce79004a2e66aff1774d595ad4c37b61d6, 224'h2aaddfe2abcbb137ebf80d35c86c7f81fc760640eec39eb3abe9ee7d},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{447, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00d5751d00e69e86302d95f3a485c357867b31c1f726021f8318330eeb, 224'h36e15c9ab9152ca24bd32edbd0de3a10e7ccb23b493c3827009798bd},  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{448, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h2d738785b04282261457a9b149a6c51c4c611f29e14113bbd2625981, 224'h6cacb7671751394b931ab86a09631ee26cd077c01af8c3491b535982},  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{449, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h121f5992ff2892a8e0b36cf4f31331fddcb9b53d1aec2c7d9cd887cb, 224'h406a219f572c58baab779d8c386fe8e84857024a21c01f949505a668},  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{450, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00c28e4e9a7f4a96f22bab95a3f564099ec46dda7ed0d1568b3474fa1f, 232'h00a7d93ad705f4604bf82dc029d2257917d1eb7e09d4799637bbc31661},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{451, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h008e5a9b74c35d07b2dc788a9baf13764bccf2570a07cb4b51e52c36f4, 224'h1ebaa0563536f7ae6337e446f9ff9940901b4b1e6c8a6af283d56b5e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{452, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00975b1ef86996b5362792d0444e1cb8c64fb583b91477853162ed7914, 232'h00abca04859e3df4308d9d40b33798c2f0907dd073ee7587646acb2f2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{453, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00dcfda67794874a4613c1597658dc52ff8504de9db45a2909894052fd, 232'h00eb8fbc6e67b20309b9c0c1315bd2883029e049b77033fdc0be6a0e89},  // lens: hash=512b(64B), x=232b(29B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{454, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00ad39c764452e94c39dc651bca149bff4e37b7e1856ab3d40625f952e, 224'h0f454f1ed191e8cedcb9c290758bd4b9747a32b814852b1da419d1b6},  // lens: hash=512b(64B), x=232b(29B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{455, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h009ff602d8037ef12b2f22858411a992a21c554fe10e07567338a03412, 232'h0092d174d805bd0eae1093b20c4b3a74f9e09dab0a292d4147173874ea},  // lens: hash=512b(64B), x=232b(29B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{456, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h5041006f1dd06d3bebcaaf4d10e1371998d871c04fe2f730b43ec025, 232'h00cd2ac83465809b3c658115d286a8a00f67db8a1068f84ecab418bb0d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{457, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h00ee587c28d2210b0cff7d47ac3509f590053320e547d3e034df9c9a50, 224'h215374b4e8541ae4974974ed7575d2c1550d924708e303c0b744ee77},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{458, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h00b66a579ea2dca40e3a48074567af7daad34fd784e3ed097d1b39569c, 232'h0094a2b72c713c109153863ebb71a8cc80f57094d811c13fa269e14a42}  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
};
`endif
