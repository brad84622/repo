`ifndef WYCHERPROOF_SECP224K1_SHA256_V1_SV
`define WYCHERPROOF_SECP224K1_SHA256_V1_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224k1_sha256_v1;

localparam int TEST_VECTORS_SECP224K1_SHA256_V1_NUM = 248;

ecdsa_vector_secp224k1_sha256_v1 test_vectors_secp224k1_sha256_v1 [] = '{
  '{1, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 224'h2ef983fa542b64472e2bc405d9eedd861acc9a7f814fad8275ce6b9a, 224'h3459ba4ab52164883bd29eb6ac7e6d22ac7d302c053dc39684928ef9, 224'h464bb0fb437b06922073e124528486e500b1394a05e86b0bf58aa70b, 232'h00f2819cdd8f311adae3930586d1fb883ae071cc8d60435904ffb9d872},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{2, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 224'h2ef983fa542b64472e2bc405d9eedd861acc9a7f814fad8275ce6b9a, 224'h3459ba4ab52164883bd29eb6ac7e6d22ac7d302c053dc39684928ef9, 232'h009868b57ff5572fd854ce7eb8b8513a1c54501e8fef97540291059a55, 232'h008ece23bafe5a9456b59d1a17a03da1dbf825cbab651ec7d143d9b70c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{3, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2ef983fa542b64472e2bc405d9eedd861acc9a7f814fad8275ce6b9a, 224'h3459ba4ab52164883bd29eb6ac7e6d22ac7d302c053dc39684928ef9, 232'h00a3588793e8c156fbfba20ee28c8dc7242460330a71868f6c68988db4, 232'h00b3db0f3fa566afb6aeea4d3ed9eb65e91b1a6bedbe77b1e27154aa2b},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{4, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 224'h2ef983fa542b64472e2bc405d9eedd861acc9a7f814fad8275ce6b9a, 224'h3459ba4ab52164883bd29eb6ac7e6d22ac7d302c053dc39684928ef9, 224'h31ec5c59558df32ce76d49cce64d63bf85ce4c28b20bc3b375fd4a9c, 232'h00adf21d877868bc754eaa1db8847caa33ddd9ace6fdcea59c1e37e32d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{5, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 224'h3fc04f62221710b2a8510cc9cdc437a622fc0dca8509d7bde7e55ce5},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{6, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 224'hc03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{7, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{83, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 240'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db00780000, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=240b(30B), s=232b(29B)
  '{86, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 240'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db00780500, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=240b(30B), s=232b(29B)
  '{102, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h261b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{103, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db00f8, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{104, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 216'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db00, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=216b(27B), s=232b(29B)
  '{105, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 216'h1b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=216b(27B), s=232b(29B)
  '{106, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 33000'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db00780000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=33000b(4125B), s=232b(29B)
  '{107, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'hff241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{109, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 248'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba55120000},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=248b(31B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 248'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba55120500},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=248b(31B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h02c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5592},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 224'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba55},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 33008'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba55120000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=33008b(4126B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 240'hff00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=240b(30B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h01241b54acec345f866a6bc2c440169db878b78d3e93e7aec93e7ab26f, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{153, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'hff241b54acec345f866a6bc2c44012e3e6d2deca34fe065be6513b4e81, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 240'h0100241b54acec345f866a6bc2c441f1a9a2922cb084b9a076ce678cf778, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=240b(30B), s=232b(29B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'hdbe4ab5313cba07995943d3bbfeb3f305a34d4463708faa83824ff88, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00dbe4ab5313cba07995943d3bbfed1c192d2135cb01f9a419aec4b17f, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{157, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'hfedbe4ab5313cba07995943d3bbfe96247874872c16c185136c1854d91, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{158, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h02241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{159, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'hfe241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 296'h020000000000000000241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=296b(37B), s=232b(29B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h01c03fb09ddde8ef4d57aef336323f822b82dcb53f10d77b25055a0709, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'hc03fb09ddde8ef4d57aef336323bc859dd03f2357af62842181aa31b, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{163, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 240'h0100c03fb09ddde8ef4d57aef336341a8e159c51d8853690432a2e6c4c12, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=240b(30B), s=232b(29B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'hff3fc04f62221710b2a8510cc9cdc25abd500fac45ba192e4c7145aaee, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'hfe3fc04f62221710b2a8510cc9cdc07dd47d234ac0ef2884dafaa5f8f7, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h02c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{167, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'hfec03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{168, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 296'h020000000000000000c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512, 232'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=296b(37B), s=232b(29B)
  '{169, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{176, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{177, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{178, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{179, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{180, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{182, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{183, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{184, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{187, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{188, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{189, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{190, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{192, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{193, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{194, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{195, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{196, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{197, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{198, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{199, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{200, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{201, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{202, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{203, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{204, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{205, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{206, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{207, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{208, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{209, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{210, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{211, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{212, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{213, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{214, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{215, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{216, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{217, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{218, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{219, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{220, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{221, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{222, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{223, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{224, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{225, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{226, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{227, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{228, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{229, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{230, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f8},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{231, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{232, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{296, 1'b1, 256'h682a0fddb418968157ce8175e0ef497ae3ead6e9dcd822590da315c7bb337f67, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00b3b20995de5790b06f1baf8aac6cb45d240b94f8386ce5cb85fd767e, 232'h00f9ed86660b3f8cab18aeaa3c7ccc171781c37849e202f91234428a67},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{297, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00d185705d14349c8135580703fa073448588c3fa6c3f4fd1d259baf0a, 232'h00f265b8ab29519fc6d01c64dd10508c25a0da8a84eba301b3a45c988f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{298, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00dcc8e76934dd8f2898ea3913dd13ff819bf11ae7ff4092ba02e5810f, 224'h2baf248326573f71cf0bee75de4bef569d993cb2fddd723a779682d9},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{299, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h7f3fe54fc07dcfef793d82276f4d65683fb2d97c0c36262880dd83ed, 232'h00f2e7f13c3cf4f08057e61d49cb1fa771c0bfba07b61a15a569e2fc54},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{300, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h3e2f81e04eb857268f9637f4c74fc186acff0caa606108abf3e589a4, 232'h00f454f0afa411cc0b6e1851c99b5569ddefe283c15911df9081527613},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{301, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h7c0828d863ce6d6913b1c286f73953e4ae012e848a052e82afda0530, 224'h0d7e7befa3c03caaad5d76afa887f1e90a46458074f3655268994f0a},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{302, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h5e0d4c378d083719d87502c5d37d173169143d3caefa1fbe9e0c0de2, 224'h6e64b7656ac29958a7ca2b83ae97504ac97b4fe7f79cbed87ee43f51},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{303, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h008b7d2b774cfff76b2af7e26442a9ae208e1dc6a34ef834f4b4457544, 224'h1277305bc63a6be1c7391843c49d84b2c09e4559915bde823ceac80d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{304, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h73097b86f4e6d993d712283efe20722179853ab4f28cac9133e12574, 232'h00b9fabcad69137c3dd65e77dcc4af68fc3962dd068d51d38fa458dcb5},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{305, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h0426536cadbf410c017fde31a0774b55f65ecaa4fba920b27a18263a, 232'h00bbfe0fadf37bc81e674d0dd585a79016425b433aa036a8bea0f0b5f7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{306, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h008118c784b1ae2bb122cc922c6d7bb12f1ee74476a337d0b928416a72, 232'h00bb6f13c2467282ff0c7b9edf55309ed4ba724465746603c295b9eca1},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{307, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h0087f59675df4fbd38e286a30a1c283d16bda45d64d59d5398050d0535, 232'h00c841b0035d9dc8a52303954b50b99451963f89944516b28cfe13a0cb},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{308, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h6d53edf91ce58bdd92e12e2d8f55d7637edd7ee59ac6e78381ebeec3, 224'h6d5a0743de3e5cad36e8894aa07a5a07a714370051b692361ad3debc},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{309, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00f1c232db08b807c9eeb2c08a9fb12cc43f501bd9307e5927ab5b868b, 232'h00b326a28d3829937393e2bd7010791bed95d84fa35119aa3a8a7e587c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{310, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h0e8620fe1b96c708db18bef7103b1c950d0b84fa50288d5f90606b5c, 232'h00cca0c85563f2a3babb22e0bb27aaf0c9bd21551d82acfaa704e60cbf},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{311, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00a0dbe08a31ec55514eb92e8812c4aadb3be44a46b70b0aa5f966e408, 232'h00ad82b9591408fb300fc55db29847b54e3501ae33709fa174e2104aed},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{312, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h675357659ae8e6b8380d4d84bf9bec14378337ea445efc5796e94c03, 232'h009804b36633faae3d5d576192904fdc24abd07bafd15a85e5299ca021},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{313, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00904ae6242505e55f365fe5616dcc0928efe3c3745487a8f066cbe59c, 232'h009e1b7b1b9a0bfc1a12c4ac979077982bba97d9d90b82be4a943187c0},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{314, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h6a9c1de2cb1969901f38ab2e521a5a4c2d054db43851f2a175f6712e, 224'h40d588366e72441ebf1b1cb2e3516dd500b3322f7ec9771c3d0eb849},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00b10e9f30ada774daed4b4ed9138f07448d1638b6b3997596031f739b, 232'h00d67d07dc32141aa5f6826d22c8a108261e52eebbc4c21e23f8e6db2b},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{316, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h5d4dbf8017a04f12d9502e63718677d241cf46cfca25413c38f38f62, 224'h077cd018618cfa428887d8cf9cc49085a7ef963b8fd01d5aaaf862a6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{317, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h1a2c2331eb8f97daf2157042ac472119bc45d661fec664483a1fc81e, 224'h305c423b008045a4f5dc1bbdd0bb7b29dcd29cd389e52a4a7ed5ac27},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{318, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h45e512bbad719cdf4023e25d5f02b9f82d3fa254c7a1389378018f95, 232'h00a9e4254c881cfd8cfd4cf8f64621a97ef349ad648f3d68b09b5fd0dc},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{319, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h4814fb555f1fa664f7c9fa3f345181866afdfe0e0826d43b63265c26, 232'h00984dde5455253c4ffb35116cada8f9e8b6f2f2dcb5e456b3fa0fa360},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{320, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00851aef44b0869b4c0f3d7d5926e6799f094ab345bc03166ba48f6aa2, 232'h00d228916088d12e4a17e499c48c0ca8feefc8b264e22122f0144e7b77},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{321, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h23bbc9d0e3178ffc71fbad8584e166aab86c498597cd1891bf407d6b, 232'h00d8b80633d631a5aa06197b14e3fc1f76778db72f721b6087a131d68b},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{322, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h593d30711700976c78bb617a2029d0b433af7b8f706856ca1248ba27, 224'h07ea97204b37184d723520069e83c27e53142a67bc9e68e777c50072},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{323, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h49285c90a8738e3092fbf78819f5b562c7da020e4881e01fd0b6824e, 224'h33044f586ac7ecdb506e1ce3f3a1abafbb44951565367c8070541369},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{324, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h7049f7f70a97bc356803cf49695b72a82b2a98b70ff1c026ff01e2d0, 232'h00f152ed9b31f1c90b06c36220d8d4a557c1b95a55b50398a47e88be8e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{325, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h1a8960b59b53ff42dc42582f58fa0d853db5022422b6885393168dff, 232'h00979477b5a23092cd7f90e48372b7efa4a78e53d1c224279b45158619},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{326, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00f0635e4b65dd762ea99b62dd8ad719d68c0ea6d5dcd02f5454735e7d, 224'h606d10db9561f5895d4ab524fb79b475580d29ecde7fdd1bb85c5b4d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{327, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h3408da6225d974875437816e5c9aa7f2dcae06b42da3d03ff92f94ce, 224'h5201beea5fdbcbfff8082937c32d95ed1a9b89121c2ed94097d73f07},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{328, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h4b375c050402389b8c7e60ff896b3ec60951b7714a7a0f89d754558f, 224'h6b1a9669881f83d75229d3cfbc4efd8d86c2d3ab2e2e8bcbcfae844c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{329, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00ac6c28591ae72d7f27282598d214a8abe7a0deceb3420f0c7e2fe7c8, 232'h009b85701bcbb2a80f72111c8ed8c182bfac5bf7816ac3e0432f2ba1b7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{330, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h2bf7cc09a7405cc9ff20028aa246322acb9d05ed979c5f67dc0522ca, 224'h64cfb2076f0773e5a0a89d81a2bac2dccf2341e0f82f8d6dd23ea425},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{331, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h009ada9fb763f99aafc2e49fa8d8d25ef9a856f9556d864ddf540e324f, 224'h7568bc71ae33acb7e200739c8c5dc622413106efd81443d7e42439a7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{332, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00cc81edd6949a519f85dccac80fbff7e9687d3b470a2680cd6f208f60, 232'h00fabc8d2ca0b84a66ac1bfc845b90c724d5e6da26c444bb3f6950c004},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{333, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h37db84341c99735661e277d8b17eca9833b253be56e22d5eb300551b, 232'h00894f213e4218e208284bb4152ef926e7b7740eac72b1816fe6ff57e2},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{334, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h008685cfc397575b4519102ad8f6e9950389a02ffc3e3b151616e6c057, 232'h00de04d0948d1e8ea4bb7ddd38c19d3a039688d9b5218768a9e717ee9c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{335, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h008b4ac0a09b785fd09f67088687f1fe7604d7e7dfea48917a6e14955c, 232'h00c08640f0386d64f18c31dc4b1a09bff70c508d05258649226b0cae71},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{336, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h6671c4f541bb626145bc2fdf8aaee83477048efa22d0bb25d3a03b8b, 232'h00c36bfe072281fdbb39ceb8899d71347acd22d63f011d29576075acb6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{337, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00a6757619dc34907429497852518eee66309a69e899678323531b037e, 224'h0168342d4a621255ec49b2e90d87ec583947afa35f04d972b81fff93},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{338, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00bdf013257440075b018e68a60a4353d017303dad825138eb8a2a58d4, 224'h4855f2391f313e7a6fb3a78f00eb48f0435d45358591e9a2bc8f5351},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{339, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h5cfdcd39f1a1cb8c259323823896c23f25d3354fdbad446d51006673, 224'h0bef5f32aa56df10f062d33b5e8408a9c1281c002c8f325242a62861},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h06b9c9328ee02d7828eb73697dd41de06619cb0581f16d6d224d0491, 224'h0431999d333bd4ee2bff37ce9094cf33e72696456122e11bff431482},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{341, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h009eedfa8555c75abdb6113c8af62ad9f501a4b0f1d302c2e2330ab80b, 232'h00fc9034a89f32a5c1e2962694981a13f11296f497a6fe6132ba710d82},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{342, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h008e7c79348b3c9cd6ed186c97d6986fa4c505a5d11e4283930fb64cf6, 224'h5be14fb89e87b3d821d8f5440b1ff7648a56fb9469ba801c5e57f854},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{343, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h30901d4b952d7c59a14a5e4c7c4c420b53295d6b9738111471103ec9, 232'h00b83f03ef8dea9060adb27de34814c12d6759a011f2bcceb5e4bf9f92},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{344, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h630e6f0a1a29e979aab89c830c4ca8cc9d848d5c4dd821e35a43aa76, 232'h00c27dc32fbd2fd6342bec1389bf63c27150f6bd72480b3f7289a1ec91},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{345, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00ebbb7fa96725acaadd8b6760fa1b66052817d5c5cce6c29cda9f360f, 224'h5a9cfecd47b0c014f6d7f8a669f409e96e4536a3600990bbcaabff77},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{346, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00ed1f449ce9fc545706d286b69ad395e9a3ce6bec58ea8cfb237b8469, 232'h00c746f27a705a8bb629f57d7417bf33aad3711ff31243ee5f91bafad7},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{347, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h009f047e69fe223049f4512516af3f40dce646763b2e02bd26ab75cb3a, 224'h56dc557edfa262734769caaa8fe27cbbe916a4c659da490df7b7e65a},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{348, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h45373e696c28f8d2e869e51c5ba9a8e76dc04015f479e49fa354b626, 224'h6a1f35a36ec1a1d032b48dc98f711d247459d9148d61a9a6a6884d0a},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{349, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h0086740c5821490591acfd5e13ffc317798fe6924c1564cee689a3a419, 232'h009a8fa36a94fbaaee93c743994dc82d58b4ee19079284cdb74fba7246},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{350, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00d6195954e66c78a0f8ff4d76b00c495eec59e693e9f6816661804d6d, 224'h19a6d0dafe4a069128d17cefc716158e02f0675c9884e50ceadfa575},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{351, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 232'h00838f95addf1212676e8fbca5cf34d525856116a2e7162658fd384446, 232'h00a4d53d1f7cdbe6d71393aed1c41c6d5aa314b553e86f8169b5a11543},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2cad534f3a9b9f7af75ef6b52b34e98b39afca1f76cdb3a3478d5e04, 224'h05f4b39f0b8e0e89e4d21c43d7046501cbc5506344f717487860c76a, 232'h00fffffffffffffffffffffffffffffffffffffffffffffffeffffe56c, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1f4},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h0626c8135926a2ebca46bdba2a88c99ddab5367f06ffe11ff9c58dac, 224'h296491e4e37f21f84e28993dd0e0896cf56fa05ed411ce670d74257c, 120'h01dce8d2ec6184caf0a972769fcc86, 120'h01dce8d2ec6184caf0a972769fcc85},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=120b(15B), s=120b(15B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e65c9ff5718ade2472f6a60a0932455772d6c6dc17a0fdb9dae48bca, 224'h29d6f9569efae6aedb8380a8bc8075b04eb4491edde3514af5bd129d, 40'h0100001a92, 224'h6b40cfab3ff22bd6ef6f2b1a28398acd590fadc0b1c3d530f69e2736},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00968402f95fd321c0cf75f78edbd2f8c836f2d8b55952b820f7a0ba34, 224'h354db2bda50b742a03d972b9063f455ab0f6cf6dab448b33f540f922, 40'h0100001a92, 224'h40e62110de4b8ede6ab17d2f8ac1bce1b3230f4bb3c676b2caa9150c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2f874521547c06dbcb5dd575632a45cbac3ccc69e59ccef1a1652afa, 232'h00f014b8c953ffd4e3f157130293b0cab1739a9542543a36e90b35177a, 8'h02, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c48a1d6cc5f68b379f875e4971723299b28089019afd67628e3a6bf7, 224'h09c63f963d2656bf864e080cda07cc5d30e8f4ac61bb6ea2d5646b0b, 8'h02, 8'h02},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00db7a161f1cf83a215b43ab283deea50bf2dabf29d38277ae826f14b4, 232'h00f6c231b0fbc035998fd72431475d0c1c7ecae43aa2366f3afdf5d50b, 8'h02, 8'h03},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b621d2678163deaa6fa425ec3f7a3936ce24bc71737bad547668c500, 232'h008a6d3abcd5c6ebdf88fb90b0ff3da086b41f2df5f33df5b50b9ae879, 8'h04, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d263f43fca0fda72b3f6bb521e1bba6d50f392b81b6eeb7312a21fbc, 232'h00e95f160949fa569352497e88c56f7232f204f1aade752d8b3f21663d, 8'h04, 8'h03},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{361, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0092064e58faac9017d5fd40dacfa4da86459156c8876780a993dc8351, 232'h00ce6a6c3786b87deba14855118156f0a9af09fe82999e81f2dd46e0b6, 8'h04, 8'h04},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{362, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008a5913b8da46091e1f3521703a129057582c16c60b781353f0c2b3c1, 224'h028c5efb2add74557d0f17df2795ee6f374482473a3b7b0904f6b147, 8'h04, 8'h05},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{363, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008a5913b8da46091e1f3521703a129057582c16c60b781353f0c2b3c1, 224'h028c5efb2add74557d0f17df2795ee6f374482473a3b7b0904f6b147, 232'h010000000000000000000000000001dce8d2ec6184caf0a971769fb1fb, 8'h05},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=8b(1B)
  '{364, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e8fd619638ec64e34ca3cd9093afc5937dd213acecc22cdd5552a1ae, 224'h6abc8dfa960b55bb3282c625367fb542ccc5e00b21879192ad1f7feb, 8'h04, 232'h010000000000000000000000000001dce8d2ec6184caf0a97176b2887e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{365, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00fd2b95781249901d53e78d7a1c18db65cfbce5e59d1e01d36fce3cbd, 232'h00976a445f957cd6aa009b052fc7bccdac1d057d35d8e6539f30c98c15, 16'h0100, 232'h00c183060c183060c183060c1830622a02a3783996c5bfff133f76b2df},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=16b(2B), s=232b(29B)
  '{366, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0092f0088eff3b24fd6cfb8d99adcbfebb873c3b15fad012214d22d64c, 224'h0b7b8a94a75b60f7bb4130ccc01297c7a250091d78df6a04c3cda624, 56'h2d9b4d347952cc, 224'h0135fa9cb663a24b634b6c650b61ea744182b35e059463d8479f4057},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{367, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c9d1d50e5a5efc6d387beb9fc7aa8a73fd7597e7f2b49c8174556239, 224'h37f6d59c22426d5d6be3c0ce305f80bb8f912faf9dfe9ad843128ba1, 104'h1033e67e37b32b445580bf4efb, 224'h19e619e619e619e619e619e619e64a257fec15d1aaf17fb5d03bfc17},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=104b(13B), s=224b(28B)
  '{368, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h41a2ea107b28cb0dab233a102ed40609a68ba7e1c1b1cd85ac880ba4, 232'h00aed24d7da7571c9d1934e11c919783872bc6cceeacae25a0bb50e2a7, 16'h0100, 232'h00bc9db5f704530ba1cc7ab8d5b5b0255d6a7115ba6cb5e94d54f0dd8d},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=16b(2B), s=232b(29B)
  '{369, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e052de3ece2d4bf492b7d5a427bcff08ab178416ffaf0706fd9eb11f, 232'h00862cc16f03150a4d90cb778f40f648398ab9763ad0fc86988e866943, 104'h062522bbd3ecbe7c39e93e7c24, 232'h00bc9db5f704530ba1cc7ab8d5b5b0255d6a7115ba6cb5e94d54f0dd8d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=232b(29B)
  '{370, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00fc64cb84f8f635864a29fec2897e8be844e54839d8f20c028b0f4ed1, 232'h00d1a9f5ebb38cfd8a9449a90a6dfbd73faf9c60a440919ab56e5dcd10, 120'h01dce8d2ec6184caf0a972769fcc0b, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b52},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=120b(15B), s=224b(28B)
  '{371, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00ca0b442aad1e1d57c43c67d7a648797f344233537b8dae6ddd248d5d, 232'h00e3994babccac8782cc18e56ce18772a2add8ec4d47fb807756390877, 72'h009c44febf31c3594d, 72'h00839ed28247c2b06b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=72b(9B), s=72b(9B)
  '{372, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00f39dc37388cb4c34fe5d5a1f2aa6041c4c108ccc13e42c61f0c418de, 232'h00adb51ba0d123842cbf2a83a8a75e2a3d2bed11adf11784d15278c550, 104'h09df8b682430beef6f5fd7c7cd, 104'h0fd0a62e13778f4222a0d61c8a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=104b(13B)
  '{373, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c8b6ea8c530305db5ad07d53d51d61858a13d2bf766541040e7acecf, 232'h00f255573d8521b52299bdcbf2ca5cdd4e00bb14dec6a07b7df5a56e41, 136'h008a598e563a89f526c32ebec8de26367a, 136'h0084f633e2042630e99dd0f1e16f7a04bf},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=136b(17B), s=136b(17B)
  '{374, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h49f6f1d2a600142eaaf7410097c1a644a91349fe8677963892d68c86, 232'h00a0dbf7abeb84ac9b5b2129b4b7e4baad0989c990321f33e5edf1ced2, 168'h00aa6eeb5823f7fa31b466bb473797f0d0314c0bdf, 168'h00e2977c479e6d25703cebbc6bd561938cc9d1bfb9},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=168b(21B), s=168b(21B)
  '{375, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h4cbacc728670e4e1df367749fce32c6a4f17bc634bc52f502d44cc95, 232'h00e0a864b52cdffddaeb70ed9f073484a45858889c58e80ec8007e9fc6, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{376, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h4cbacc728670e4e1df367749fce32c6a4f17bc634bc52f502d44cc95, 232'h00e0a864b52cdffddaeb70ed9f073484a45858889c58e80ec8007e9fc6, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{377, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h4b9c0cf9f218f64d1317ffc18caf11797cbb431550816b42e658da6c, 224'h5051333576ab8be2753bcfbad797b29c0b8eb76b4b310bb24f3c6ec7, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h74d89d2b42107a17e0df7430a84102f0c3befe18e59ea9ed5aef3195},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{378, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008981be0db57c743232f8a5d30b419840c4d38087d66c501597f737ac, 232'h00b07a341cac19c626da4adb9f3119cb4439e954b1718a7eae45f7a933, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h2a179e7ed670727c33ba8da63fe226140a7fcf62d2cfaea7ea59d1d4},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{379, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h69f46cfddcec6520e4e65590c64466c19cff0f581e13ed401d4f3470, 232'h00cfb829ac4e52055461d0785876d78e3d5889a7749be663a6bf08459b, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h6d50b1cb505189520a6901a895ea13458ff5076156c27efc00639c35},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{380, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0086ae72267749417993992aa8724e9d760dc3962b2ad01ebc28019fa0, 224'h5a107cf5332ff42f5516451f2298a362a894d95ba849d48ed389ffd5, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h0f59ae2e4259dbe0997caabcdb25bdbe8d6df67f433a4651342d5219},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{381, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d39979285ed39d2250c5125305868dbd4274b8a603d571e3537c2ea5, 232'h00f7c67e822535efc4c1021b6b312c34e4d60be2e89984e95f5dddb7de, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h5e10dd8d9f91876988f21a2bc2fefa4df57ab4efc82ca41a773ae802},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{382, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h5329099622fe9e1008c891fff3ba768c6d764d420509fd232830603b, 224'h2d9d32aff3af504eb4389dc7bde4f9c4c5fdac7bff001d6da369104c, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h511eb0edc14410a1c38d655e04e0c99cd8af84d8caa0ffd69da2dc44},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{383, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0090d1161f4794186cc6d0baeaa03f63e84ae61b3428712cd561978ecd, 232'h00acd7e006ada0004b6ea0f27da9ea26791a94292e57e3584af0de87c5, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h11577274428aaa4ac5d23552e64d35c2e45667773fe77fba629f873f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{384, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h326aa12c68fd569b573884a97b899c197c18fb9c509782be8b18011f, 232'h0082d76e993348dd4de2440a6d7bbfcd7461729a6ac70a3fade02fbd8b, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h2fb159d4c8769a346ee620bb1e5027f2aa0fd3b1d8b3a2411c9b9ca0},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{385, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h0633d37de65ad8897f863b485babc75cb14175692597db295e4d2beb, 224'h649f25584f8f9f3121549431e1e3ea5290ed186d443ac4b53df57b14, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h59d3622af6be99859f0aea85aa20e669ec373992af2856f37dea777f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{386, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0093f80c5d235dbb8efb8622bf70716316b021ece8a37d2ff33a422cbd, 232'h00b0fe70e8e87e04736a54a943d524b3ef27628d7f7688e901fdb25f40, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h3296bcaf337a66617b38e2ab65833612cd0bae1b7b3e670863dac215},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{387, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h6bd84040f3c08088a7dab45cb4a455a8b5336a00f2b2899779adc048, 232'h00cf5d1bdbb1042789adeb363dbd7c4f776560f7d3c6ff24e58d0709c0, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h1b468ea6fa697becc552ec879c3e9ffdd72969403d5fb745bbd7f366},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{388, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h6a942adc74e5a542beb5a9ed73166bba16a621fde05fad8feb93041a, 232'h00b9d8e5797a2e237b2785c36f24156dd40d3ed35064f8878bb6db114a, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h244b2ee0f3acf3ca0d086215fbc12728516ffc93c03d27a601d31a8a},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{389, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h74897882013164324092db05bb1d2e0d44386fea0ad1b2eefec19565, 224'h0f28f541785399eb1b825131e82b18da9a30049686fd4af36fff43ce, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h5625c3f523582b7986ad997a8488acfbfc4b2db75913a1fa4b437ec5},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{390, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0081a4a2c2c959ba5ef743d32f173b1e24567ea1c37fc5cf6e36b02577, 224'h079d37fa3c2f8540bed4d6465ff45ed71878ba86cee8ffb4776231ad, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h148bd1fd5c6502009ef1febb26c374cacd3a62e7f3f232e21f145115},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{391, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h009473345d373f2e5511b33bdb3dd2335c0eb3979eeb8176972ca6312b, 232'h00940b9640487c1b5c0c501c91bbebf037e42f43970ff57b55cf8d4a7c, 232'h008000000000000000000000000000ee74697630c2657854b8bb4fd8fb, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b52},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{392, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e34c5ec17254bffb619c695ef1f57b337307178260de9e3afd1b0056, 232'h00c45191abe124ff2b7e7444e3e4828bb501978c4de01d9570d6758e77, 232'h008000000000000000000000000000ee74697630c2657854b8bb4fd8fe, 232'h008000000000000000000000000000ee74697630c2657854b8bb4fd8fb},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{393, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c1ff9c2ed13e9898adce894b574a9c1a07507e90613001e50a787a04, 224'h578ecd045261a7121e12ce909fd2509ec3cb2aa9082e7b80cc075f44, 232'h008000000000000000000000000000ee74697630c2657854b8bb4fd8fe, 232'h008000000000000000000000000000ee74697630c2657854b8bb4fd8fc},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{394, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c8185e31d2c92b095a0bfbaa54341919719c17694fb4189277b8c203, 224'h01d456a7ff02096789fd426737f735b050a1a6c918b3a0cf6cf0f838, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b4e, 232'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86564e19100f4833fd},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{395, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h20683d2970e76ede44f92ece6a6c2ec0a165724ac3bd725f968fe039, 224'h53baf1f5521c63bb4b938019f6b82625312c40a247cd92561114e886, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b4e, 232'h00894b5a17a0c6db3c25793c14d7be760ba56af3833f9339d2ddf72ff1},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{396, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c73ef8ec74b35b83942ec13f90b838147e31e00c84c82166fbee4a8e, 224'h2adf5032da443a8ec22a4cff4c3a4724a79ace6394048237b5bd6890, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b4e, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b4e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{397, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h342a7eab53183ab55771a1dc973d9514a475546ee0f58f10251d4ce7, 224'h55116ba58412a175c71122063c4bf6d774adb1d2f27ab3b160d22b32, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b4e, 232'h00aaaaaaaaaaaaaaaaaaaaaaaaaaabe89b3748410331f5c64ba46a76a9},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{398, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h6e812955a9eeeea8ebeffff30463446bb4bba9f54687be4a7cd7ad31, 224'h32c67a10c00f31e826e3b8bf50da9826bd4aa29270c004f4d5c5692d, 40'h0100001a90, 232'h00d23c374d75130c4148d796a3b817b58f9bc8bb03b5bf962b2ca2a1fc},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{399, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h14d87a664bac68655b1767aec2bb50c920f92c31eb07d4f08cefd2b2, 224'h618d1fbfff7dfa24e85b3ac5de8e433618fe56480698113a76915f80, 40'h0100001a90, 224'h050bc5eda83286e4e8506020be6a8eb2d500ea3be9104339e91396fc},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{400, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h1c04f658b6f346d883578f43b7a7022595805df36ec9135fa60ff384, 232'h008b3363c603485d2c56ed870277319d18426c26fd600306f41fa64bc4, 40'h0100001a90, 232'h00e14150ae375f5c042821b2b1bc3806fe885461d0cadd0fecef622e2d},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{401, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h29e8873e1492e132461dd827cb9d6bb0b824789ef3d5c7211015f0e7, 232'h00ad90890e2805e13c5fb2968a5770cd580d6d13f8dbd182b8e8c2ade7, 40'h0100001a90, 232'h00947e3ca712b14ca9894b5a17a0c7efddeaff84f1461aa0419ca1d30a},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{402, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h1a7aa4f0d18ca3d2b63b70f8045fa368c08dc9ded1f1a27ce43aa052, 224'h4923a32e3a6627159ec389f5adb1aa4bf1c8196125ab5de07db13050, 40'h0100001a90, 232'h00e3ca712b14ca9894b5a17a0c6db56ab329525d6aeb501e2699a4957f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{403, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h31158fad37ccb15efd5002f7b0aed5c56f31c099b6957fd1a6afe0a5, 224'h19d786ee55ca132dbf1ead663df5bf62b810ed324bc07ed9dd5c9ea4, 40'h0100001a90, 232'h00c794e256299531296b42f418db68f87d7fb859510baf92dbbca97907},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{404, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d67cb3bb26f994c8a6e591b821245f5e118b2667b7f75c9251eef200, 224'h61b5696a63106e89fd531b9ccdfae032a668fe274bc1cbf5be1bc200, 40'h0100001a90, 224'h12b14ca9894b5a17a0c6db3c25795ee7825cdea7d37ffcbbcc8b03df},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{405, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h22b01f7ed9019b0d96aff38822cf9cd7644ee1ad0cc5d1b2a3f67bc2, 224'h16b5dcda155b053a914f59cf86b39e2d6882ba4757a8ca9d84b88d66, 40'h0100001a90, 232'h0087a0a17317277df51e86bc3a0bfd4a589d51772d3e55d7ef1cfa0650},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{406, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h04f39a7ded5b62d429e3af6d2718457ffd87a9d00f4b5389e0230848, 224'h57b0cbadb8326c12a2fc15a42206d515011ec6e5272583e5d2036c1e, 40'h0100001a90, 224'h2dc3c8b28aecf3beb728695c47ea27593723a6811531134649fd0ffb},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{407, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008278a0f8fb890f0df8c4c72c40d55cb5ff8c5c39f280c917b76fa5c3, 232'h00e4e68e0b21853347f458409c88cd160990486cdf2e0d094c1c7484d5, 40'h0100001a90, 232'h00c4a5ad0bd0636d9e12bc9e0a6be0297a3c2baa840541f1a22a4b70f4},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{408, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0080a9a9352af442fcfecb93e8566d34e455b0bffe53b30ddc59a7f10f, 224'h33291dc141ceb06597ef3e091dcd75413484eea32aff99af5d2c78cc, 40'h0100001a90, 232'h00f0a0a8571bafae021410d958de1cf1f3ada061aacae6dcaf3300f012},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{409, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a824ae928cb209d3d4143a8cd10a7b29d863150a5482f873972e6031, 224'h12f9d12f2fff94f4e0a5b9e3e5a88bc21b2d09da15584ca655c31094, 40'h0100001a90, 32'h55555e30},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=32b(4B)
  '{410, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00fc53f6e5bef640cdfb14fdfe17172145b795b6daea5d3eb94a995c82, 224'h353627058219defd06caceed9b10520ac8e6a06ed793273c585a3ab6, 40'h0100001a90, 232'h00b64b7ce572ee917838a4cd1441ce7a5870cb872b6e1afa7d474581ad},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{411, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h5e423679db282576cec351f1500a4ee1a3e6bc146b76c147c3798fe3, 232'h00ed029bdb0474eddaad50e2a6f2780ff184b33f4c38c03738ed6c1ba7, 40'h0100001a90, 224'h39232f26cb0fcd6b2eeb69ba41b9ef00813616da98cd16e2ef21123f},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=40b(5B), s=224b(28B)
  '{412, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h038925a04a7e62c3f709ae4150051692290405fc3e2c0ec2eb0de428, 232'h008d7148d65237c36fe18e125447adf9189793b86f5256e915c52d44d9, 40'h0100001a90, 224'h121c0384a8d015f000000000000021bc8ed98db7f846a8b77b820ac0},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=40b(5B), s=224b(28B)
  '{413, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b5ed1385fd9206c7e5f60ceba655e8f0fe5f46cd058ea5c756ec4296, 232'h00bd7fd5bd557d4fda0853583b5ab5aae1b5fc2adbecb9c0a8f4e4ad55, 40'h0100001a90, 232'h00c0384a8d015f000000000000000166177c01689b50dc2ea136641829},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{414, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00cf7680caf9081bbcf6ab137781f38cad821115358a9f14d20e343a1f, 224'h500dff2e5067de9fa32331bdad78809dd195dba19f9157fb0eaf4e08, 40'h0100001a90, 232'h008070951a02be0000000000000000ef4625166fb1d6c7b3d0f6287e5b},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{415, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00830814c8b60123572cf9e740f12de791198bc9be1f9439eff154e0a9, 232'h008e098f637ccfc6687f95b54f08cf9dbe246cd0b638a938d545a3df91, 40'h0100001a90, 232'h00a8d015f0000000000000000000013a7c7074b3a182ae23e0218e57a4},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{416, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00976242536e189112598b48a6cd3603aea2e573f95f780c04e55ecbde, 232'h00cc06c81713c45020788448e707fed861bc6ca97d8790a3ca93fc14e2, 40'h0100001a90, 232'h010000000000000000000000000001dce8d2ec6184caf0a9716866ccef},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{417, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h1f087f752f3e023f66d5487d9123375d11161b516174455bcc18764d, 232'h00ba3f6edb1ffc8c5cdb338bdfde9363361db29df1662d375959260a02, 40'h0100001a90, 232'h010000000000000000000000000001dce8d2ec6184caf0a971214a53c7},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{418, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e4220766ddba093f8d7b44b4a2c6631808e31a30eb019a1b50d94ee2, 232'h00faecc0a837e7e88a96f9848ec32bb52032fb66f1aa171c3fe7819f52, 40'h0100001a90, 232'h010000000000000000000000000001dce8d2ec6184caf0a970f69fa4af},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=40b(5B), s=232b(29B)
  '{419, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h1fd75eec503aa7f892d5133b8348e1888a40f1af64aefa0b480010af, 224'h76509a2b5607ee7a1d87cfd6f9e8cc5255b783809e56ddaa8f4151f6, 40'h0100001a90, 232'h009c9197936587e6b59775b4dd20dde5f4aa113c2fb1dee02a32e0621b},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=232b(29B)
  '{420, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00dcdfd288cd39527cae16e666d7c1ab01fd548599251e9c7dfd3195f8, 224'h1e72a8cf308f14ac7cff3eeb189e29e56be9cc4dace858299d2a6ab9, 232'h00c294f85b63b7c629862a1d3afbf880caf92695bc763a51bf8b3450ee, 224'h17dffe0d34cffc00054c58130dd5bd8e069e95fc4acab8bccdacdfe6},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{421, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00dcdfd288cd39527cae16e666d7c1ab01fd548599251e9c7dfd3195f8, 232'h00e18d5730cf70eb538300c114e761d61a941633b25317a7d562d57ab4, 232'h00c294f85b63b7c629862a1d3afbf880caf92695bc763a51bf8b3450ee, 224'h17dffe0d34cffc00054c58130dd5bd8e069e95fc4acab8bccdacdfe6},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{422, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h5126d8509cc88bd0ae29c97062b8ba4b416906294a9331bc678dd362, 224'h65171023f5de2d1c8a2da0080f50b29972875fc7c1bf9428d95aa704, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b52, 224'h33333333333333333333333333339294f6fc1380f5635516b1532397},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{423, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00ad0435d05538bdea3b6f75bd2157af6e581ba0470e6b176fe48fc43a, 224'h45e9de57c4f65768602c6dbc3f48232a3ab5d8a475509a63727a08ac, 232'h0086c0deb56aeb9712390999a0232b9bf596b9639fa1ce8cf426749e60, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b52},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{424, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h721c01fa7cfe06059affd4de9c75c7b556cf7f02490cfc4644b48b1e, 232'h0093db5689ff2282693dd1e19ac2fae301b0d410e5b8ce778485216545, 232'h0086c0deb56aeb9712390999a0232b9bf596b9639fa1ce8cf426749e60, 232'h00b6db6db6db6db6db6db6db6db6dcc25d28f1fc836c62c22c794d7f1e},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{425, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c8ea63c6afe1c64474e13b6d579fd9edf20f75b9ecb60150c4041ad6, 232'h00adfa14549ecae5920029195e4c5426038ba70058c7f3fdd394d932de, 232'h0086c0deb56aeb9712390999a0232b9bf596b9639fa1ce8cf426749e60, 232'h00ccccccccccccccccccccccccccce4a53dbf04e03d58d545ac54c8e5f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{426, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h7f6ccdfc4bc1a0a699d938b6bcbbc7930b1374772c64e458a3396105, 232'h00e1b8048589069de732a8935f3c40e1dfb9b215ef95ae173eda60f03c, 232'h0086c0deb56aeb9712390999a0232b9bf596b9639fa1ce8cf426749e60, 224'h33333333333333333333333333339294f6fc1380f5635516b1532398},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{427, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h060a436d62c31fe65f90eb80347182d818c898155f1c821c829a2eaa, 224'h45db9ff41a6f5e6a6c7ae4eb7ae1bcb53db9c95768e907c8b4d446e7, 232'h0086c0deb56aeb9712390999a0232b9bf596b9639fa1ce8cf426749e60, 224'h49249249249249249249249249251a8ba9fa65015e8de744fd5232d9},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{428, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00dbabab2e4f527a54179119636e0cbfe1ff47898d711054e668530c28, 224'h1127e0ee1ccc776155d9e957f5cf8a14f138b47c51b3b98b3a52b658, 232'h0086c0deb56aeb9712390999a0232b9bf596b9639fa1ce8cf426749e60, 224'h0eb10e5ab95e2e3a079268cf3a6524239ef04127208663a54968804f},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{429, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00ff74391905cadc0cd906fa519a873b04d46fb0a5950a6d2739b7c238, 224'h6124bc5f2538b2195a99ff9bebf89e49cf890d22096e0c9e9f455651, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b52},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{430, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00bc641827b39c4035b146fbba8c0b8b4d160781ef18ff59b4e9a0e8fd, 224'h7e772274ea9aa156c6891f4132c009191f881e6fc534bbd222481b11, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 232'h00b6db6db6db6db6db6db6db6db6dcc25d28f1fc836c62c22c794d7f1e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{431, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2e7cb47b3bf0bd2f1708f89161b9310f6b72db0245bb4bfb9a175ecf, 224'h23bbb92cd72771d510e6ffe99f40079d38b37aa1ba08db2f9e96fa6b, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 232'h00ccccccccccccccccccccccccccce4a53dbf04e03d58d545ac54c8e5f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{432, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h1bc33add16c9f6d80dbe98dd620408976c497b2bba6bb1a390c52190, 224'h74821a06d64f86ee2b0888efb032c9731367898eb398836e5fbeb5bb, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 224'h33333333333333333333333333339294f6fc1380f5635516b1532398},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{433, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00ea602b888ac8095114fbb0bfd56d2df146df5a5d664370e33b0c9e9f, 232'h00cab9b3aff24ac5b4282a7f1e32a375991028bd5fe3a8a1d211928506, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 224'h49249249249249249249249249251a8ba9fa65015e8de744fd5232d9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{434, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0083e6196134f944eb73a0239b6eb32249eefb5bc91a135e46efb97a95, 232'h00bed598f10b7a81ca181366fc087eaf48bcf47ad8ecaf720f7f72d992, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 224'h0eb10e5ab95e2e3a079268cf3a6524239ef04127208663a54968804f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{435, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 224'h7e089fed7fba344282cafbd6f7e319f7c0b0bd59e2ca4bdb556d61a5, 232'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86564e19100f4833fd, 224'h24924924924924924924924924928d45d4fd3280af46f3a27ea9196c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{436, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 224'h7e089fed7fba344282cafbd6f7e319f7c0b0bd59e2ca4bdb556d61a5, 232'h00894b5a17a0c6db3c25793c14d7be760ba56af3833f9339d2ddf72ff1, 224'h24924924924924924924924924928d45d4fd3280af46f3a27ea9196c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{437, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 232'h0081f760128045cbbd7d350429081ce6083f4f42a61d35b423aa9283c8, 232'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86564e19100f4833fd, 224'h24924924924924924924924924928d45d4fd3280af46f3a27ea9196c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{438, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a1455b334df099df30fc28a169a467e9e47075a90f7e650eb6b7a45c, 232'h0081f760128045cbbd7d350429081ce6083f4f42a61d35b423aa9283c8, 232'h00894b5a17a0c6db3c25793c14d7be760ba56af3833f9339d2ddf72ff1, 224'h24924924924924924924924924928d45d4fd3280af46f3a27ea9196c}  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224K1_SHA256_V1_SV
