`ifndef WYCHERPROOF_SECP224R1_SHA512_SV
`define WYCHERPROOF_SECP224R1_SHA512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp224r1_sha512;

localparam int TEST_VECTORS_SECP224R1_SHA512_NUM = 322;

ecdsa_vector_secp224r1_sha512 test_vectors_secp224r1_sha512 [] = '{
  '{1, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'h394766fb67a65fe0af6c154f7cbd285ea180b4c6150cdafafb0f6f0f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{2, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'hc6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{3, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{93, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab0000, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=240b(30B), s=232b(29B)
  '{94, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 248'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e0000},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=248b(31B)
  '{98, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab0500, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=240b(30B), s=232b(29B)
  '{99, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 248'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e0500},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=248b(31B)
  '{114, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 0, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=0b(0B), s=232b(29B)
  '{115, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=0b(0B)
  '{118, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b1c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{119, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h02c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{120, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf922b, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{121, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbbae},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{122, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=216b(27B), s=232b(29B)
  '{123, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'h1c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=216b(27B), s=232b(29B)
  '{124, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{125, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{126, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 240'hff00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=240b(30B)
  '{129, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{130, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{131, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h01691c723dd6a7f5d11b8c8e8bd08173428bc48a2c3f031caaec3bbce8, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{132, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff691c723dd6a7f5d11b8c8e8bd08345fcca52a9b01748ca203383686e, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{133, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h96e38dc229580a2ee47371742f7da36054f46611d4da0c9a70206d55, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{134, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0096e38dc229580a2ee47371742f7cba0335ad564fe8b735dfcc7c9792, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{135, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hfe96e38dc229580a2ee47371742f7e8cbd743b75d3c0fce35513c44318, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{136, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h01691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{137, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0096e38dc229580a2ee47371742f7da36054f46611d4da0c9a70206d55, 232'h00c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{138, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h01c6b899049859a01f5093eab0834104e71ff12bb612ad778fbda8e56b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{139, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'hc6b899049859a01f5093eab08342d7a15e7f4b39eaf3250504f090f1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{140, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'hff394766fb67a65fe0af6c154f7cbe11bbc0c7c488012fb1b59eb344d2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{141, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'hfe394766fb67a65fe0af6c154f7cbefb18e00ed449ed52887042571a95},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{142, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 232'h01c6b899049859a01f5093eab08341ee443f383b77fed04e4a614cbb2e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{143, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h691c723dd6a7f5d11b8c8e8bd0825c9fab0b99ee2b25f3658fdf92ab, 224'h394766fb67a65fe0af6c154f7cbe11bbc0c7c488012fb1b59eb344d2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{144, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{148, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{149, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{150, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{151, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{154, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{158, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{159, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{160, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{161, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{164, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{168, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{169, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{170, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{171, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{174, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{175, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{176, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{177, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{178, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{179, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{180, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{181, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{184, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{185, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{186, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{187, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{188, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{189, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{190, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{191, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{194, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{195, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{196, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{197, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{198, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{199, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{200, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{201, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{204, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{205, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{206, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{207, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{208, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{209, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{210, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{211, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{214, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{215, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{216, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{217, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{218, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{219, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{220, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{221, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{230, 1'b1, 512'hf582f7e1597d4966b5873f6fb0211f38c289b14924aa3830aa767732dbda99f309d9c9561dcb6255ac12355838d8587b8bb0d09d5f693189904337c73ee68378, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 224'h221a25eb9cc8dd66fdf156b2f6ab601ab6d9c509247f8de5d2671a96},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{231, 1'b1, 512'h0000000001b99889c891f2468c618149cb6865b933cca31eddb353de09746b540616ba69c5f5ff992c6d6177427daf1cb46a4c5c08625263a615fbf3eeaae178, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3b3008ed596b7fa276498def40d96b1eb2ffb731a44050ffb732e4e6, 224'h6dbb08c56db737e9392ff4f3a54d8b806d70af226ecf413b3465de55},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{232, 1'b1, 512'h7800000000c52e48c315d5276f18d994c345b5805aa02872c29105d1bf75f152042a782853b4a3850822714434fefe3db00a19bc7eb84029869a7c1dca47ce71, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d1fe269c3061e4b94604e8d612d70887068cc7d5232cd5a9b72923a1, 224'h3c1cbc027d33fb2451d52dce3a828a8c7ecc490a28a94e5e5bb2c4d7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{233, 1'b1, 512'had9a00000000987c9531c475b0236659fdd3dd795473bafb8f0753bcaa4bea4e6418f79cba317764c48fdfd9461986dcf668f250be9ed2b7b75afaac70ccf0ec, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h04586134cc679295dd93499311c4a8af37cb94dadbae18d8ee279b9b, 232'h00bf9170a1b65b665664cf567d40a995ce252a23d6a9f962b05e364486},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{234, 1'b1, 512'hb3284200000000930b8b98132341f68419e3262a7f2b8d60cfee7e1e364b36ed4f000bd5fcde187cde7397820b85a174025e4d54d70cbaa80d160fc9cc72d56d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c1f51009b935b4773374364ec3eed72a24b70926e0349c77862f3475, 224'h46df3d98f104ba6602f8041a5bf5495fb240e103d1bd17f2fa878923},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{235, 1'b1, 512'h3bf2ef06000000009638300311c31a5caa29197ef0d079767e66e50824e8d41e5a36f593539a6c0ce102a92493c18061c70eefb94903831d9b8ed3291d1b9829, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e822242872f1ecf338a4f773df87b67e9b21bb283acac7d66b26551e, 232'h0094d4e0fc3c6359994a6eaedddd1533f490f72ef85139f8d3b39cf07b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{236, 1'b1, 512'hef200f1a5400000000399e032faaf4b3c32d804555abf20471a3a18dc46f3917eb9072220b5d5f994d27b221346631c47eb579d69cc5e438b7e7b963bca9d84f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7fd45528eb7bfc3710e273c4468f0b50ebf93f94cd0e7a602a4929a6, 224'h46613dd1ffd85df8d71f3498001721fda4982c27a1c291359b05b1b8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{237, 1'b1, 512'h7f12580858d000000000055d6877381f726e0a9237d1c012c9840b5b3fbeb6f43027bba37a94ba5fc0dbab436b88d4a7cde6aac151b06214a00cd8fe5f0bdef8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h36d137b69171a486933b50138d1db1842724766afd25c85b0032daf5, 232'h008e700de21f2fc350a34c7cc19054cf371ecab6f7331ccecf68fca0f4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{238, 1'b1, 512'h6b4185d1e7382000000000c86f684e5386df6f2e7e1dab4d1be30ccac1ea33d4e82d455b12857120cfb411b75c8df08758216dcb774dedf1438bd137f831b27d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00da3b436908f5a82f26bc17a8577ad2a782946e3a7587b01d253b1dd0, 232'h00a6544e38f24e8117370c049b5d1f6712ea14337a94511224df4496a3},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{239, 1'b1, 512'hd40c1a66696b7a6500000000ebb22b0b1f80b394770ad61c5c42ff0584ed4c84a3d185d3c07725f0d3080b451dad86945cc9b0801c01e0b6b8739ff8ec36df22, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4314a2bd139d47be3d9fd9ebdd72a06a220219c7596b944178ee6f5f, 224'h0e6f1d2f57c699654e9c705d7b8fa3c1ccb0f939f6368bed246b2e10},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{240, 1'b1, 512'h68481d736990000f3d000000001bc2164f3bf7a43f3c7f23a875b84fcc1d1395c9bc3eec02e9aa7d38f4462d5734ca53f0db4e46498d1b8c9f9f4c92f4fc0532, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6a25643464682679d84970c603927f4a8ca83e7ef9715dd1ed84c28f, 232'h00932b78d165c225a5253e6201c0b1ded0898ba24de44b23233eb78054},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{241, 1'b1, 512'hcf9bb31b573fa12e7e51000000004b37d8761e5d50f214b30bc2b134bc7e0e30653b8debc737a21392357313d13e08eecfdefd8d37bec92b680a84f5430fb57c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h476aaa58677d9e60477cffd026c43248e2cf3cc21e8fdccb75ceefad, 224'h7799fc7af8f9b929203faf899bb5ca1aecf2492555157282dfde790d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{242, 1'b1, 512'ha678a93e12f88e59d6307e00000000bcef462484d98a07578e5106f6b5e6cd1618aa82e3797b4bf519cdc4704616039255cb3f05fc8b93e4a48e2c4cd5333450, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h63a98614a1421e2ebb278de53b61618bafc757122647affd358c667a, 232'h008edba806e0a7e438ca35f98405a8ad2d5c3e8cc2d5c4384233aef0a5},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{243, 1'b1, 512'haed2cc5334773206d7170bca0000000081dafcdf0acf2107d7c016b54b1c0ef3663c5ba78277a328ae547ffdf6ef2e385a374d9355022f24dd05ff9b357e5039, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00880b5238a014f8b44655b83c175880eb1e8307899a824ea3e07dbd6d, 232'h00a4724c8649fd74e5bc8d7fe6a9067a1376fb8e08dbdaed68980b0f50},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{244, 1'b1, 512'hfeac570e6cd1481ff79f34cccc00000000eb127fae412cf598abaa6550b4f5f2e1537dd5c5d6c57b0b52c103ec0340c9e292d0a263d74e44301efe65d505ff9d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f8743588234634dd9891f4f2f40f4e46b77f97b82dc5dbe234aa6b5d, 232'h0080656e5262bc25e158f3b78f51ae0d6a41cc8cca1aa457221b2eb7fb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{245, 1'b1, 512'hbacfc820b1f513e6a157534762b6000000008ba56a4c814c4c12a828e658c8f7d0453900871cece52dca13f4f1df23685d1bd43488e2acdda903b2e0f72b9d64, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2a2357e3d8fe34434582be4dabd58b77b388d1d52adcc664f45dece4, 232'h0094be3a369b7c2788df4587ec5bd4163c4cbc40b77de1a85e8bcfb251},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{246, 1'b1, 512'hf9f58ffc6e2662f4992e06774f928d0000000084b7ca7f7b6fb750919f466be3366746484849f67645a424ce6009fc560031052d0775f47984d3a4727776b916, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b6b0c0aba6c611300ecad8816242c415f183a2bd4d46cd7769033d9b, 224'h7750b24be02f22dc0b656fe4af377413f9453dff99226915dbb6e08f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{247, 1'b1, 512'h5f6f67fd931001c593ff6f8e5ea8faac00000000ecb4ce9ec81a128cb55bba07a9b186b28f7e787f7bfb7ea32d9047b830a99f2ac4144ee3f6e07ddf00e68646, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a5c1a75c2779f3eb83a65e295927cce4288e9d5c2132a4c7ca92526e, 224'h10fe30f0be33a785385137b57d806140a402b9bd3c1df1b57de6da63},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{248, 1'b1, 512'hdcc948cfcd6f3cd3760d678a643ab0ff010000000095bdd5dd5c0b9579c7c6b0f3e921033117737e31acf8ab117b62ee54a25abdba306c71bb0c3d60097a332c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b92b5521d1a7abe77e8524dbd3001121cf83c08017e3917bc58b5d1c, 224'h224b113779017f6a522171edf930f1b5d4f5e7dedc6d2d514fd7883c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{249, 1'b1, 512'hdfc50d9e551fd99c3ceeeadef83e2fab3f96000000003206a5e2b462805d83d6ef6280540f3bfbb229421d6f5f2794f117259f9dace4f82dd57889a74a0fcce9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ebd3ecf3aa64cdcdd171585a141a4a673a8d5de0ca087dfcdf62432e, 232'h00e0f1a0f7b8f5ac4a42632f87156ad1094079393b03f2051a9fd60249},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{250, 1'b1, 512'he4edde495afeff435a69e94a6493e4ec2c0b1b000000004c8e512f917698225b0189f732d3deb6d8c1c39b6b59e0701bd7f7605a521891358603454d151d8e7d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6c3854297e1f267b64a28e0cd6148e0fadcf85bc8d5c23947543bcb8, 232'h00aa0594ee11312f5d4767d296e5ca83df68072811f81a8d27e178ca5d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{251, 1'b1, 512'hdf8f102f7c54ce2cb6ca609ce724818f7621cdc600000000c69bb15b7c33f6b27c75a153b581d47b99de18ccc8105fc3bb697f180112706c5ebfd6fc6c8a6322, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h785ac8c956d7797ae67498775b3c446c41735eb15f3430b49f6a09f2, 224'h5710879ab83994e809c8d2cbd6f2ac5c205b4b8d6226e98be03e7967},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{252, 1'b1, 512'h3e526c3c1f02aa2e007cecd9e02f7dc3d06f361a0c00000000f8e183a89a7218d8183a928d91c6bba47d950bf841396e5fedf9d87f66671deb8d2ebf63e39751, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f1f3d016693125ba73981c8f9a1748e5dce1d9634355f26fa536190e, 232'h00b574e97def60dcd0e9177106483791b2edb4ab0342b9f5ebb957d5b0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{253, 1'b1, 512'h7a750c1372a8d9b00991182aa031522b94a1a7f4509a00000000baafee68e65ef0a94f7983cfeb9241e0b7d8fd590a0d55b16041eaaabc38e982aaaaf6eb75e6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e64f3371522cb1a5f0d1511b152b20e01deca0b3284786853cac279a, 232'h00c9a2e5f4ffde22b9d4ed0179ce74fff408ea918dda7685c7980ae61a},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{254, 1'b1, 512'hb8df763eea0cf11e9945dc5667b0147cf8684d618abe1200000000917eeb543a4dddd7217ba71e998bb9c5fd62b57509b7cdb489bc3b64f66a70e4b5c12ffd2e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1f99dd6ef72feeeda6c123baa4fabb126d7dedb64130fae3f4230797, 232'h00e441ec51dca6271b043e95753c4043d7cb4e76fdc13d6aea45fbf243},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{255, 1'b1, 512'h88670299bf6b255d331cd40c7154c438fab9fdd2b4319e440000000057a51b1cdea2812fd594a8cdd56b4f5cb069625524bd53a5f304653824d4afbf9bc58d02, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008637a09627c52766bf96f0b6cea6f2ac3eb303001c5f6fe6d628e4ba, 224'h10b66c599455d40077bb865ed43e2c2cc403473baa6d63b16be48c84},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{256, 1'b1, 512'h295422dc27dfac13c79d2028d3daed64c1dcaad525dbbf14a9000000003667b1baf41fd9137fa0bd8c3851590b206aefb6cde62fb4ecc23ae308e540e83a7f09, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h52a010a23e4f9ebb459bbe9f3057e6c19761fb99d25c9b16b8f007d8, 224'h526dc1f34444de00447ba23c76950f2c159579d548b6335d127ea321},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{257, 1'b1, 512'h118422376e38638a08705cddcdd319e26fc8a2e6d4a4d1400fb70000000005687b339ec07f51592f6e254c9b7291fa2d0302df9fb2702857e3f69bd4fba01654, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fc49caaada528f3357e5a264f2e7f970ca1b15ca5fee28741d1202ac, 224'h175e884d10d0bfd20b39311ce2c53083da167d1f3dfeb990e59ed628},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{258, 1'b1, 512'h5a4801a1f7ef2afbf8e0e76cbd6e07212568cb47638e22e55f8e6c000000003a2aff81ce04258211030942fca855cbc0ef482027b17a7ee523b15483afd91355, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d95d539a85c9edacd4e02ede27b0e0b737099612d166c637c83a9f34, 224'h59936a2b90b7f3f3da83f64dec8e347a3bfa57baadf9acea18c071d8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{259, 1'b1, 512'h057d7524efbce651b92e0a70e4454156e7cd4b696c197c6a064032c100000000768565d4af2019fe3247dba91948292af777f107fdc9c3b47659eaeab26ead77, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1895e65593d71e5635cce022dda19bd155bb9a7f2e307e5ce9127ade, 224'h121b487c320c544dcdd471d46fcde2ce5dc9d17fda70544c4eab50a2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{260, 1'b1, 512'h31ccd924b687a2a6b70f4888ea911ea38a686e56e5540ea692ca3174bb00000000246ac69c46506bd8fe924eec33b33ebc9f508d4251c459fdcee3b4c84d4ea3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b5f4c85b13b51a5da81a236f1105937f3d98856d2aeb57101b6b499c, 224'h3be74ae770fa6467f76a742eb9e504a815a4a60e74b38bcaa89f9b06},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{261, 1'b1, 512'hc7b70cc4a55d55342487a4469ad2243ef6d6b69f11604b8c12baa03dd3e10000000014df0db29a9d4d54b26f4047f3e0c739f7a260768b20589254e1235fc590, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h07a57197667a0c40423d4811ff96384c9330467e8a28eaa4c0d519f4, 224'h011062c8694494baaed24ff610e1e4227efb59a163c33fafd40100f9},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{262, 1'b1, 512'h1634df8a3271a99f360e3bbdcf789d24bf4bb03e3114ee9f0fa930541f1ae0000000008d976fb74f27eb316ce3a24d92a53833e600c353300f5c4fec6b28c581, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'h7f718615ba1d0a9d27a8c5a678a6225ffe1233ed8b417c9343b310, 232'h00cf6a87e4496725c6a2612f4034ddf4b31c7435e2fc3a163e92d463ba},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=216b(27B), s=232b(29B)
  '{263, 1'b1, 512'h8f90b6a8ecbb870dc24832b1f4719aae2d8eedd7faf97848b08d2b528abf5f44000000008877a6157344e6a9dc43b90c8e2dd7ab9bdc5237c912e094660d0878, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ba8f95a4363c493a9f78bb61dbefaa9587d028bb8344420de2b0cf21, 232'h00b3798c2d6e27a2591c2edc18320b78bf11df194b11b3fb498c595232},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{264, 1'b1, 512'hc0891fc626ef4b106fc00f5c067253f26a2868d09aa2ce029466f353ba525e757100000000a3cee37421995445fae741697659a406394c870d8bdda130080d15, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h596b74077801db2e889d3b2aaa3990fe180abc152d48528385ca955d, 224'h38bffd416f779843fad389750003eb0708112a4834c554f476a3e0d1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{265, 1'b1, 512'h76527097fb3945436a30cca60392c170abb7ddf6ddae93e3ff7651d468eb3e14865700000000bd314c31706f8e4d1d853b151f5afe680e13cf2f255b2bb697bb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008547f62967523a06c9690e5ff66c3f2254cda28f09ffccc222433d39, 224'h3d9ebf664ee551bb7b33157d6c6c5fd456bda3d4ae460215ec1a5f94},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{266, 1'b1, 512'h41d43cb27d4db522756dd682826eee8d0f60163c7f3ce67a39d89d7d89e24818c354ef00000000cab56830cd18f7bb9a7d1b2440fde06ce647518fada2dc988a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0090ee3fab9c6ce373a1b35fc135fe878280ee25e58a4bd7529e91b4f0, 224'h6451e7526505b44e88472b46eda3fd2679824dcdfc445e67f35ea382},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{267, 1'b1, 512'hd34ac40ed5ab79a4e5ac1e4081e0e47e4fdedac1555b01ab62a13ac0ae9dbc3c23f799510000000010116f328ad1db0cd68cd1db9e1b34b5a52ebe9b8e372b78, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0a530530b6a9238d2d1a3cf468986c87f3b208f61ea0486d53140c17, 224'h5f027a73f31a5cc2bee81ff0019477c542fd782ecde0e551fcd37e93},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{268, 1'b1, 512'h8b5db6db13b1f5e609965dc38215d14ccddf66a9d86505a67cca37f13cc420803c1df80f4700000000b044bda09a83e4331aaff90c4faceea315e467f5fd91d4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00beab4abd23df5e2acfff07c82e245dfa7d587d0238c2c9ab9c88a96a, 232'h0098c6507635536840edf604f9baae6408ce4d3fbee694db3abd825011},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{269, 1'b1, 512'hc771e022bc376ffbe1f513bcff11884e790e53878c197014931f6360c517ce8de1c059d091cf000000003c560cc443a6f005ea58917a52ca9bf60163afb16ce8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ec8c36335cb98fa07b983c35b7fc256f44a5aa192d6087595145a15, 232'h00c32b7a47ac6271f4593562bbbf91f9e07395a5e4d46970495cf29f05},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{270, 1'b1, 512'hd9cb55a3f1ec161bf6caf0452bd6d6c876b35dd1000eefe18378afaef6280348fd799e624e573a00000000085b3b24635f5c10770090ea935f198728655e236d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bd635a741f1f2a1d9ac1698baf5cfc491d5e3f8e15f1cacbe4ffe4dc, 224'h4bb606cf7cc11d0d7d96b83966f42276095ccc445882ed5afddabf1e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{271, 1'b1, 512'h0caacc1f43ee27ec7ad5269155a66172ac310d4e202a9b7d3defcfb07ea8da85415ac2b116e665830000000009887d6c7da6cda824528345e14a6675de23988a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00812c08622c0a09d949b7628585c4f4f2db4c5591b5da148ff46d5cd4, 224'h2104f9bc9d0079acb3077d2db58f388119500c5322cb9b5389b5c5d7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{272, 1'b1, 512'h5d761de2a231df86c0fdd90da20e5811f7bd9bebb3f1966359b8fdf554f79f0bdd32ca06410e70e61100000000ed3d4140a60908e85f7fcbd26dc792bedacbfa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fa4e1c8b0006f269c855eb495fa3a113f643fa8b1fef2b08ab145994, 232'h00fe85b8b522c7f9e8943e0f62643395bd1fcdabc892c315d108b75f65},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{273, 1'b1, 512'h78adfad2734b7baf32f4e0201bd6c3e9f6c1763cbe35858a0f56466db34dd98a0fbf5b2a71afbcdeebd400000000d3da1a5035406b39aa13c126a3946b6c6a5e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008c1d9b7911bacb6b4a09582648b992d46a1832eb006178c0c77fcb10, 232'h00becbe12b99f243766da5bdad07461b9226a8298672b4f1adb35357ef},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{274, 1'b1, 512'hf1d6ef224f72b83a109944afbfb34ae1f70d6e50eee54a91faf8ba0fc062563113d988f2b826c055ecc61e00000000554878a7e761e75fdf1ed2ad2d138b2974, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h78850a40530aa258e478e7c547d3a5e4944d3524f1676443e4dfb37d, 224'h687058e1ca478f52a30c9a3f8e2eea9d8c40599cd47ef66b9430d17d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{275, 1'b1, 512'hb33f308c5b107050cb2e513fabf8b896e52c85852fbe32308bee8b8661121bdac78f52f924cf3d5690ac92d5000000004f0f619e72ec1464166078ba3f508a66, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h066e7268a6abefe1b4b916ca51c3e958e40dc78c3661313e0ed2e77d, 224'h6404d8a332a837f2ab6bd13e3ee4aad1e9307d449e7f9b7d6332030c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{276, 1'b1, 512'h0392f8c2dc961605c5693d9452731b6a8292ff57d6995aeca0dad3117459668ec7809dc09cf154170fcd624be50000000026e3d92dfdf1a2abd09392468117c9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4eca73709a67c41603ca5af494c8132483ffc2e0bf171b52de5a5e81, 224'h2c79137cd2add3ce3a76792270e347221a3ad786eafc2682b39bcf95},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{277, 1'b1, 512'h9dda0539bfe47c75bc00b014dc6046c9db5d7a5723acddaccaf2aac7a9250b732a80cd948409f132d1dd65cfe91600000000d53c76be9f75fc6927f818acdaf7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0178512f8844984222393a63263e0a009601869e632f07eb7470aa05, 232'h00e32657cded1122cee0a4f66ff50a32da1f05de4c5e217acdf5eb6fe2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{278, 1'b1, 512'h572e1d736d78c42eed5ffabdfb25b5c7908aa60728ddb3d36a24c285db9ab996433827aca9e23716c3baabbbb4527600000000b9c1a728fdb6f65c10935e9514, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e2c7bf1222ca23a56492873c2d3fa6c7030cc166d693142dcea272b6, 224'h715a4c82fda4404217dea6c0bbf3ac24f8faa2b435fbc6d51a32c4a8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{279, 1'b1, 512'h81b675425e8c528a0a51b23413c8b796411a01b207e0bafc5bd2a46b05237be84abdae1ebd492fca053bf7e3133392720000000086ce63108f1dc5a3b34c575d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h49886a8c26c91d649cbfecda6ce8d1441e764c66f5d81dceedb6c5ba, 224'h4370d8bcd4f052fac9491d62850b6a6a85d5acc44d9248c3dff30bf2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{280, 1'b1, 512'h11c203ef3c8978266a73147233f7c9c9d16108a07847ff587f1e865f28519e7a161664edb56d9e791fba0717124717b3c90000000013c59e26ab63c4a99b871c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e1ae225e1aeca40747ff3e7ad1f75eb9bc90d637160a7f58ce12e591, 232'h00b97cbea3a9323110315760b7e2ede496514b30f0eec521ffeb07a634},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{281, 1'b1, 512'h5de83c97136ff31a90ea5053ff256d522819626ae3734c460ea7681fbd0a94538ed840f3bfbf8055756e761d8149786b8cb000000000f37f36e4d32d46cb9bd1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008a93b87b46512544fb9a7af5c41e3aa72e40235ef87ccb7108daae48, 224'h157db617ac697df407af7a11626c52a1af7ef189514da39918c43010},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{282, 1'b1, 512'h4a5e1e8c073ecb2832fe0d0df42a72ce225ea97ce093ed320aaba00cab25ec3e90a6aefaae72ad40273d7309e40582f40a37c1000000000b1e8576da0eda555b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ebdebe6388b9f460fce6d84faa67ded1e864ef09e77ea3ce58a5deff, 232'h00be5052033eb40380c2b1325fe97dcc55841e147a89f02a296b4505ef},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{283, 1'b1, 512'h9f920bb92b4527d54ff6877b80c81585dc4d3d1e96fce780b030f9f371f8a1b68e2e7a86536acc3ce96737bd5fba0ff669f6b1600000000000b5868a36cfe6c5, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e85d0667972d003c82afb9e18b702357119b4f38401a5ebdfcbea88c, 232'h00eb7b3e5268a4ce6280f72d7e9a3d74e5cac50b1c3a5296cdb5a49d82},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{284, 1'b1, 512'h99f941e73ab790b224ce0a799133f6b04eb9bcfb2fd0ec84b8e7d5dca6ca50d2b1ae4d31c57e2e54f97f59b6a10d0758cfb3e46500000000909d4fabd9d1962a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3d243581c0874fd4eb4d80f896c5067429ad455314881951ab5ec6e3, 224'h0ec47aba08ccba88c1a6ddc289f595bda08dc2dd34d12dcefb68094d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{285, 1'b1, 512'h202e258cee0bca789ccd4c29f3835362b6f1f53faded0f1d58f4ff768f6202a6de3ee3b922546127fecfdf1c0446605751df9b7fbb000000001a8a11a3e383f3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h75c966bbdcef9157d47a134231229f9f5ee8ce458775fc747d4509bd, 232'h00e344fa716e2088d95a55d02a978a416da10f22a5cccf35a2863227cf},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{286, 1'b1, 512'h8c4a184638926ecd8f6ae279181f9171181295757e3eae5b5a0de2fc0281358973a355e4820da4ce0c69db549c72ea007f80ae990565000000009e51983c039c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00cfdf599e986d770b73784d97149f9945fd16d22c302bb796156e7fb4, 232'h00c6409785047b0083f008771b40db8502583208b61c8984671acb0929},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{287, 1'b1, 512'h92eabef5ab4296dba863345a2f11c2bc8d32bc02731323a19a88897aa1421f384448516975b6397a8e627fd3cb5a5dd6ee3c50226b18860000000077b18d5c83, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c53c4aeec8f2e7a5cc0e885a6031aa1a6c1b7b7fec83b5084cbe291f, 232'h00b0e6d10a8fd86f958c3b0f4662ed8ca0d6eadbc892aac4200fcf8315},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{288, 1'b1, 512'h4cb05f07197bd719557dcfbe1edff395550b275100cb073ecb4a0987621f83a5f041996f63fececb77a30cccc5f8067e36f650f7defb611b000000006a949e2d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2386550d6e75350bcc32507bfc9beb9c26d72ff82f671c1f5282e98b, 232'h00a55b8de808c4359fb529b80a80d9fc6eddb5ce08082c3b677c689991},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{289, 1'b1, 512'he744eaf4e9c4c17549ca3907721df98de95b69d07d56eef509d4740a3cb142bc61b6c4d108676526d5a77188977d924dc9a8adf6c01adc35d6000000007f3077, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1fbd192d955ce02b64a3be5bb21bef22b53a6c6f9576d8f889b09e4e, 232'h00f5a9b673a4ee5aabf1ca8e8289f25b62a3e08b956f7418c03e2d3031},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{290, 1'b1, 512'h4fbf285c9be6083627ef151df0d2c5fb00b6edcfc44216a30467a4fe268214ab66dd9be898bea57b48f6499d09d4beddb7c9e8bd813fe7c1cacb0000000054f2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b80ffba451db9fc2194e450bdd43bc0f53a7d0f4a78900c09fb8d9bc, 224'h0124eeeab9035b6c845959e70b04d1e187d554807d6751afabcc1802},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{291, 1'b1, 512'he698cebca57a541614e179f28ba51cf82fa0fb4300f81df5fe22b635eb4441b496a36ad280999f503edded3ae1cab1700758b5ae80ce33dbf25c7300000000e9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h187fb026ade3ad16dd4b2813e8ebda433cb6cc3af1615bedf486a9e2, 224'h6fbee53fa884d296f34f7719f74919434d1b7090c485eeed2fb8fd6c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{292, 1'b1, 512'h43f5ecee4c9b5bcf2497d9753beb1eca8a01c143f8b50518e83bc7f3f62d049b03430a6dbc9236d54b7ef5475a232e3de9160e9649e3c8f46d2f1f7900000000, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e598a16fe12da79e9814f6985c9a9334010f287dc9e38de857ca5fc0, 224'h19e0ed54f0e08ad091a163b4c7b86d0634da2c86a7a8991f5d8706d8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{293, 1'b1, 512'hffffffff4fbe152fff953f198736b155220dfe633b6fc7aa5bb392cb96cde9fc658b17828d0d04ece0f6e35ed6bbf357b86665cac7735a3b9c85c038d4a85019, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b31a10480e397c8aa46f52a0f2fb5c22ebc0534fba156718b50cf6ea, 224'h602004df4b47a2065130ca3b05f1eb02d0b37b79b04b1eb799408346},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{294, 1'b1, 512'h47ffffffffa19c2322e79638701c393ec0df74b5d27fb9ea7cc3e3dc8badffcac83dd8c409a22c2d7a64b5693f153f60264487aabe5df546115cf2eaae415ac0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bc47e242d19dcc6321913980d73923e430bc6623d219529d586619b6, 232'h0081397dd2f52811b534ed754a937d904f04a7de278fa3bc8926de6946},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{295, 1'b1, 512'h391dffffffff5a981c0576acae266e7b35ecdfeddfeb6db903e9f4eab200dba039b146517f0c5b418d096addeab6d0962a6f77c2a2a552748b788c07796553e5, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5be0e0dfb26b1caa88f866504aa8e76f035a82abe00028d962bcfafa, 224'h3c3c1df06026123471bed324ca79c51b28b3d10b1ce877cef21b852d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{296, 1'b1, 512'h8c8ed3ffffffffd5bc0cf4859c831b89860c28ba17ff5a259b6982325be66498c4ac3119da331db0976678878c73473aec528a7107d0d9b1a17dacb9a9237b1f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fe79d0cfe455724792cb5ab0580ad4f2918c1403ec12f0bdd2ce6528, 232'h00f1357cd4afc402994ab868b0163f41701e0f00e561fdd97e0db6f7b9},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{297, 1'b1, 512'h531341a3ffffffff263c81971e877fd7cd8308b0d536d7fa3c88e3beaad332ef664f76387e4c43dee6c0a06423b18d1b1772f65acb4f9b672b97a648cdd25929, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1858c5d857124cd703e7c2f5e99d5025d6d979539c6f50b1d00fbd34, 232'h00d94a5adb6d9c5001162620415541d49334fb929bc86a350ca4591195},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{298, 1'b1, 512'h2639a8ec01ffffffffb54d98af88ba2ae383d69bee2f5fadda599d58796fc766130e3fb8f4ec1afceb8a1c1faa3ad305a0fdd65796adf8ac579c1306d5f0195d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e6b2ec967cfa25f57234b9ef1d87c5945502cbbd5831c862f00774d1, 232'h00caea26368bffc8e562b2bd03aa6c9dc41c529659fefe6597fce9cd9c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{299, 1'b1, 512'hd9753a5a8b1dffffffffcac9aa24c9d687a2088ed837789e72d457d0bc67f54860087c3f0509744e0b461f88893e2de6c757705670006c9e9e8c4c3757fcb160, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a59b438b2472074a93a289b33f5b13e604977dd3ab4d744d08e1061b, 224'h699574a17dc8c7298c9321ca78552e5128ea801d056f387ba42f7a09},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{300, 1'b1, 512'h9a6bf9edc61a22ffffffff703f4706318ef947658ec44c90cc1630c916924f1635efd88bcb900db41dad160ea33f8176397bb8593e19199207ca7d57bbd28305, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h748481709c6882c4a130193834a57f4bc714906211ec6cc12c400dff, 232'h00eec6c9d5a06786f821a8117eec3dc025ed3ac74e39e98a16a4aa285c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{301, 1'b1, 512'h4c18a4947b15af08ffffffffb9de1de3873b4c26280b1286a51715dcfd1242208ad49b2aad0864d5a4529e4a653d7a6355b7c1747fa9d876159d43806661395e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bc8991b506997403e123136a9c140a4336364733b0815f40d1dbd5fe, 232'h00819503ea3b4c07fc157f948f6949705d560a881fc1c6af4b7391765c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{302, 1'b1, 512'h6e50953fea8dfead2fffffffff824e02147d010595358c98ec376055cb9ddc1dfe6d3874cf38e8a98ef0664fd3b10605bc14506eb7e46460c9db81b10e2f6730, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1caece75c8e31bb0c5cceb0842f23683b8557a97036574ea88ceeabd, 224'h645ad3276aaee22b693647f00dce5f91a03b678b789b667cd3b8e751},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{303, 1'b1, 512'h1539fd34220ed16ae0b8ffffffff88a04bebde47a3a94f1b86bc687c2ce7648caa7d42ac8693b5704e401b7c9f4864bbafe3bcf761d862739eaee02516a0d707, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3a7d582068aaecaba945203bc445b3312e5cb40886522987aced68d0, 224'h39b3c612b6743a13bb2ffb83514d690cfcb9a7055e3a993cb0863938},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{304, 1'b1, 512'h69e3c78c7125bdee7184d6ffffffff274929ae7dcfc4692b84880a518de1790a758005ef7d4e29377cd891eb08e9fda55ac99a11b4dc9a15ceaf8887ae941fd7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f773c49fd0645716d16e559e22c39101df266cdfa7cb61ce46f85280, 232'h00df6109fd77a241031cf03b376e001d8a3cd2a6b646edbf9e578133f1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{305, 1'b1, 512'hc3b630a45b21b937bf78ef4affffffffad33da42317364a1090ed4446da7738caefc807ed99c92f85a6f6ba946f99284d4b9793896bc5e0b6f93cf1b09b35a6d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h79cf893f66f7faa5ca08553ea03456107e7bb391a5e51260cedaea84, 224'h32e8e3509468da7216c59975d4f3d5493848a03f864b2332044e68d1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{306, 1'b1, 512'h14f3b0fc1795c9d400d904ea0affffffffeabaaa40c2f532e33f6c61620d23188712a838f9bd1502b2a5c321117ed6007ccb48b375c581fadf340b0d7edcac93, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h025ecd1a7ab765fbfd25a6d7cd3c461e17f465e6958bce9f492b7a5a, 232'h00a1ca95038603d302761e416935acbd6b716a316c9b79c57d4053cb79},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{307, 1'b1, 512'h386b3f08bc91c7e18354f3d46de4ffffffffbf492f2bf174abad52337a99f29dda6891d96f85efb667480bcad7d2482ef7f32a314b4dd39576ef560bf01fefa0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3d14a4c21ba4dbd338fdd8b15fcdd0a9228f157cfaf2b09dd4f2aa67, 232'h00e1640e8bd2a6110dc18d6f290b7325814710c0dc88b76f127c5e9e21},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{308, 1'b1, 512'hcd86d593a60faa34608d5bcdb2e878fffffffff06003c116f812eecd35fc6f3cccc1dee24c5cb89cfe9d41b0defa4e5d16b1d9aa4897e6efc838a8a6dd5f22aa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h258dce916ef78b9d8a87beaf6edd35bcccc08c5de488586e1b7b749a, 224'h4ff500db4d665c7062179c099b2985a814f99fbfa44a3a709024d589},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{309, 1'b1, 512'h7939a3e06bee091634b535adc98afd56ffffffffeb0206c5b2cf892d2c8fbb5a2e105567cdc4447b476525488611a085b870e498a13b891cfb9a66ad725273af, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00cecf0aec5357749f357c459575298a3384dc4ac381438ff99acd9993, 232'h00da7adb092a6890e0918c235a62d4a949b0cae5e57856975108fb2b91},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{310, 1'b1, 512'h180c134c29d50916f2c3b32bf43382eeb0ffffffff6178b5edf0856813b75ccbb537c57758d3e55c190bd8e648a79c5bc6a62e45f2f037aeace1733bb7260707, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d77f2e547fd68d5db314901da1ff7ecaf3d0c17ec047a974a7cec33e, 224'h443a97afdf882272bf0233c8c4a8d23c9352ad89b1770c26240f6650},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{311, 1'b1, 512'hf2694ba9c9a0d83faff7ff2f06f0495682e8ffffffff1d5cf19e626efbbb1425dd286e93044edf262236a46a82638145b4d15c18aa6e1edc919e22bff3a9c5aa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d5dcf93e6e1b93323ea2642d3405a7423cb04f59c03420193f394886, 232'h00ddd5842e4928ee4b5d77d43d4a4bfc7f991c899727b75fc941b52995},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{312, 1'b1, 512'haa2db4394e6e52a9f0485ea08186ed648a109affffffff19fae34ae6524a6abf956c07617b15896bd3dff11cdaed4f9a2769cb4dad0b0e007b66c06fda3f256b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a9bc3ebc6ee34421326711ce29518d02bd403ead806a3e4502efa0ce, 224'h12610b89a61689a8eb6e062d2524278155fe499ffecc0e0d940d48a7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{313, 1'b1, 512'h59ce78a87d80e90e1e6b70def3179e12e78cd5f0ffffffff11eee1f43a7030f096c301beb60d1fc2be04d27aaec7c385fb9aadcd6fa37cbea40783569080dffd, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c703c508784ef71b596dcd61c5b01b45c6c69d2b36a5a3b7701e5976, 232'h00f05444a777204118f3ac2afc92d0212831bf7002158e7c656f4c07db},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{314, 1'b1, 512'h5d07345f237708f45b49a7286977f331a27c8cc58bffffffff492a29a714f16596215046376e8d35cebaaa06b73f14ec0731a0607ab89c4edee5ad7f575c93af, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0080674b740b64d383677c049a6f4baeb214f4a6b5933033853e634578, 232'h009b3a804c75ed790e31966bc25730b7428af8c73c65fb503c06c597eb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{315, 1'b1, 512'ha6d55690f7fe8dc6a67ac00e5f136dab1f6855b53643ffffffff2585eedbf8e7c3db326f7fed8c48851376d7b1a34dfd79aa6837d19b05becbe8b8d122d1baf7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7ed658c30f4a0dcc894c39f9320f59a185509ffee45eac6023577c7c, 224'h47ac94a501806d5adffea9fcf3ccd8cf79f3cc47eca9fe38fc4886b4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{316, 1'b1, 512'hd42f5eb7f42a9dd25a5d9513de8b6ccd5bbbd029263799ffffffff3baff5bcc111d8fb4f14fc4aac37a1dc5633df840644aeb69aa87f390c090e6730bade402c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h397f669cc399a91da96c16efd233f6fe60d1b7caa397cc257843b30b, 232'h00f19375fe66eae4738ec9dc5b7ef51cb33d4cb258f36944d37dd245cb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{317, 1'b1, 512'hbf0fafaf135ee4e03b991ef87e6e9377150ae255e043de57ffffffff10002deb92f4bf4c1770933d3137b0165ebcf81c8c3387c21457e0fe0c39c7c7947837b9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h537ec369b3f0d891e166f6c74e5d73dd2c4822210c5fe5f978c34072, 224'h0b183c48b5f6e69245cb76e1e2c39663eedfb74ba9538739ac495ff5},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{318, 1'b1, 512'he0dff3b5ebca4c971f1da5a6726d24519e4ca71f45a548d85fffffffff415d9ea4bcfbe4749c275d6594e8ca8b76166fc90eaf2d9f466b0f0a5ed8c14eef030b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d0ed7159cc3a79988f3c279287ca8ed10bb8f02c8b5a6204aead1223, 224'h75ee1e5c00e81899bfa8545edcc64fdf707dae1f61d976d2f0883777},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{319, 1'b1, 512'hd9a9dae1785ef8a49d7c81b0637471693412a29484ea1cc780d5ffffffffb70ab50279ba56f6576dd87ea0cc08ed51afd395238936b4aef7284700c8d5aa9f05, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00cf43329a9781db8044a920758e58399866fe7748c0f5d6a3bcdcbcbd, 232'h00d9740d2dd716290ad4160345bcd4af03af01c44b610b1e5953199075},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{320, 1'b1, 512'h75c7b98cfddf04426dda027ad897cd5ba9d5318c27288ec0f6fb67ffffffffb744ccbcda470681f3689c70425ce514d035e05dd133da5c2a104980f4ffb91014, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ab2e92c8c9143f9d8da3bdb1d935cce3ab60ae99b3ccfe863b15d14, 232'h0088c89302e8a9c591c6ed16b1ae46f966004d0b2685449842e291d742},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{321, 1'b1, 512'hccfcfe85e6d12e377ff1bec515ce149719d86cf3591b3dd8d4344022ffffffff60380790c2be6a944f31e63ee7b421a42ec5ab43f84f05aadc5ae5c42a6455b9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h04f60f8450b448198cf7981116de06d4c4888cd26be3a5947092238f, 232'h00cb23fcb33c14f089c2ae030146d68fa65eb9b086fa792f95be8ecf35},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{322, 1'b1, 512'hc445da85686a33c8af5997da14f197df87bc3ff9f277b46831c87f8147ffffffff0970446a79a2c801e1a6f9c03509ae9b782a31b3b15dec03f5789a8345e14a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f270f7a70a96a0f916c7530c6dea7178e6c087ddbcc60aacd8a7c553, 232'h008b2c378554121365a180ad4edf1a12e566ba55eeabf525356783e603},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{323, 1'b1, 512'h6a94c0cd0809f1ee1c23039f735f24a0a006a0504c295289507a9dc93e34ffffffffd7127f6a21cd1ec975e05b1a8d78144da6293f4440723e7d6062dae06a1b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0085ad01b236ca4a5451969242e16165d322428235a2af8fdcd6c4c7b9, 232'h008eb2998c5e0aaf279793caff59a266ca2068d94ebf77bae81fd0fb6a},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{324, 1'b1, 512'h31599cefc10a3c6d549bab5b19bb49d01fad30283d27c8a4905d18cf61e045fffffffff3efa7e2362af0fc827c4bf245dcd58374b350097d26ac996598012290, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00cffdb8d64b5b84b490ff73d77e51cc7797bf67c5ee0a4999def17230, 224'h3baf4b34e1a35e9606a460b395063a554264a9c43cc302ab5abf473e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{325, 1'b1, 512'hefe7f8f35a94b65eb3a9299658db8b8256f29f2df969035fe5769c11e85c9b7bffffffff61e57fc3e05c9a1eaf760ce1b13dc6ddc5516048677e1fcd420a6427, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h66cda58a5a6ddb9476e36dbad5df542be88d7e447bdc3dfe1d9e8b2c, 224'h0d99d387486a964ebab4e29bad583e46a5a200391d1065768a4e35fd},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 512'hc5c3daa9bce3e7422af1de2fdc992b34f5c8ef3fd448b45f2426e1677feaa86aa3ffffffff6e9d87ba471035c9beb5d2c94f3bb0dfb4c48298a8615840c621a6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3200761902825bd353908accd2be6b482645646971f96dc490706a37, 224'h3ed77899efdbe418370fa7998df3b7c924bed6864535277f805c894f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{327, 1'b1, 512'he36dcaffe4916e59e41b560c2961fba82290150d1b262323c674311ef6c87564c8aaffffffff573ce47a2b2f25bd4f6468ef2788ede75cd3b7293ad2bdb46617, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ba0eff0ee46aa9fca5ab8ad64aee4037931d3ad0b953d404ef9f7bdc, 232'h00afdf21df0dcbe39c2f5fa9ef7e1a2bca87d1213d1eca438929ad8982},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{328, 1'b1, 512'h3f4f00f697d80c258cbcaaeea0f4fa499e0675441a078d32627378ae08c27dc9e8b60bffffffff59976ce86a303743b716e53422d7a17166a185fac1b7722d2f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a20c6883fc6ec1ca4bb378ac88ed670a742a6284113d5fa3182a1858, 232'h00e0a73b913b94163175d264224cc70736f2fb8e8d58e914b18c921323},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{329, 1'b1, 512'h21b10973b98ea1dfd2b0d7bfe4adf9d4e8616759177daeef38d7aef0d95d226ec8e1da39ffffffff43f8e40342757a93e72541afd7a58ea2205891c13c72a8e4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f2f4af956b0c5409949d377e9bc68e4f1abef7969b518f8beacf27db, 232'h00df3a7b5993d2393ade70a2cfc1e8671a78ca4fecb56425a661a2d2fc},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{330, 1'b1, 512'h3be3c1c0f8b8f6b9c476455ceee9edbf99283f1eab4a28ace9494eae8da166e4aa1d5def8affffffff3d69a06db8c19c0984bdd10df6ede19e4214183d3b0762, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h331a1a553494f8524adb4e8a722d558965fb703ae432bf3cbdb255c2, 224'h5ab6e3dee6a2516fc4e0ac88e6dfc81d2bc37c98949cc03e521d389d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{331, 1'b1, 512'h14a2049293367e5ace79214bfae58e1007b4977ba9dbd787dd703160651e580fc6de8759ef1affffffff483224ed924c7a2906cccf6b3b39e1af044f2a7047fa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00867135558e06e19796ebce8e3555c607a6607d46f7c8da6b8552ffc1, 232'h008e827e8b9a4f74efeec7d7ba5c23428fde0227df55a1efc179a353b1},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{332, 1'b1, 512'h745beae01e0b877f882a42a6339b12080d956dfd5fa03fc87f6c99096ae69833fab59c416b092afffffffff5deea8d387d1ecabbcedd6c2334cf7eaa7aa55d84, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6746903ca095bfd3f6378a70092723483ca190b2392d8b1ad337969f, 232'h00f33bfae0835c23a80ec9f33ce9a9035c192836a0b2fadd347d803f96},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{333, 1'b1, 512'hc09dc1025bb9bfa3ef093eb420b7712374f3164db871d4cb44b8ebbeec2d5b415a73427419c5e399ffffffffb45643293f60ae63fb9ff87c56cb45252c8c7c29, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7fc0d8739ecfe349e506e71203a6e60e628a1bb0c67d5e574cb8831c, 232'h00cf8bb1557152c57550a0fde6571456fa752782f7f92f7bb235dde39f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{334, 1'b1, 512'h5f9b29b201a8f63acd7387dd71844b5ee67ca50c5a76a2b273a80d167abbdb6727992779f49b848976fffffffff2d0eab3e1c8f8be0d76338c7e8c92174b32c9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b4486e3139e0b1542892db3d3f51b0524894e19cb00cd07b03ee9c97, 232'h00ad9728d77a8b7b4fa435b3345847860c332d65d8152aa6503ab18755},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{335, 1'b1, 512'ha76f6918ab70eb9171fdaecc8add5917f130dafbb7077543007be1aa2cd3e446114f1fed5989c6275e0fffffffffd7f5a47bd23e9cd47f4572a1d1146b38972f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00afbbdc8e50e801ecbd2e3705079717f4f9d69f3b3d85215aeecb4fbc, 232'h00eceadd4e2cc9cea10b56d16a03fa551fec3eb808bd8d9f0926d14ed3},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{336, 1'b1, 512'h1694c34168745c74ab9fe8224e6058e045c73458f7e43e3884e3ed466f716a7406be99e0ef57710a1cac21ffffffffd497d0337e572f1afbc8b6b4f41a873e22, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4a762f7d146f9eafff5ad11a6978260c818b801c3488dd60411f5cf6, 232'h009ea77512585620ef2cfae8b8c9d8171229a32197e1949561bb75a049},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{337, 1'b1, 512'h3c28cf3e9527af87b483e6261fe32cee8e67cbc04b983566b27f8419a932186bce21c021eb58c8ecb0b707d9ffffffff035e36909fbfd832447041be74d2ab4d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h227fe52b579833feee16c287d29273e2256df68aff0b94d2752d877b, 232'h00bd79935e5faa8e9356622fea0135ecf796daf60333d5ab125f71e512},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{338, 1'b1, 512'hea6682cf1dadc5f218d6530a15452aaee8857a4318ef3da3cab58358a2e5d0f8fde22dc704453fb8056d224426ffffffff4335e1ab7e6e6c5f3b0a789528694e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00cd5365983eb165db39ba0c66c3a45b2ce1370c9ad14a9aa76dd4633a, 232'h00a8c77ce42ab1c888a6b5d04b71139fd882328622e15e80252e5cf7da},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{339, 1'b1, 512'h0477828c9cc5710ded82ab21dfa5887f29edfb47548a5a99ff8315da76be5f67922c0a5de1cb7448a3a79b214889ffffffff7dc823ffb5d2fbcda33e63489df0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h54d6d44373f7dfc98455a22cd39a0b320fabc33215216b37365b5a16, 224'h29cc690f2467c02e07bc416ad47204975af8c5c3346973f2b03ded3d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 512'h17dfd1c9bfab4afc7d5ac126157041f4c4ca4a04aaf17c45e47857c384fb415e4362041ec3e91609325b7e4c9fb1a3ffffffff9d3efaa9406e392a0dea1ea309, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2f5048c9ef9f30da7cb3fe4624552200f9e57a46d79db0484a0d9cf2, 224'h06dad3a4682725852869a1a459bec865661e1a38a9e546eeaac7cb84},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{341, 1'b1, 512'he2fc500440f25769bdfcc82cca36025aa6e5335d8653935dee2cc2a8e8a37c8a886885663c7da8224d2e807f62e1f039ffffffff2aa58c5c932713706022af2a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00abbf0a02332fbea779899d31d3abd2d22c9c02d4058ced639bf06c45, 232'h00cce0570f3812e5cfcb23376c554c7fc35dbcfeb623a7958c664ac6a4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{342, 1'b1, 512'ha5ce1cdebbed43dea085a592a1ef6c0881660e99434c6f3d6ec24874bb6cc9d56400958f7f95fdc15d3dcc870056263b85ffffffff9f3ace8f83061d0410f802, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1c30cb8bc21087b77eb1216ee8629e3676d925f1ae15077cc631da4f, 232'h00ee998157bdefb77d1044e983a6afec7d91a23d95c937fc5c6548c989},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{343, 1'b1, 512'h6ea638f8043673b9b6a79ff39b5d311774de5f4d697e5251ede52feecabba85d705f25c58b7c2efc844ce598d1428d22e4b3ffffffffc75b0ecb7283d80278f0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h43ee11a7ab62e2125e765c2ce5d4f84704183539810512268d87f195, 224'h65897e54025777659ee802b39c6bfd5ccc5706a9d1b38f95c078abaf},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{344, 1'b1, 512'h7cd22c5fec3646707603f858ccd785676b3284b63652913e5581a60e0c262034285489fb945534b7f2578b3e64e7b956bb6586ffffffffc05edada940cffb928, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a1fe3f4d3f43aaa3dcafa79ed99fbc045c11c352caacd89f0f63847e, 232'h00ca2e37bd2c13b9fb3f8a55b7a67eb034240395abd39fecde75141336},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{345, 1'b1, 512'hd289f68304c484efc5008425cbf00039a52c7b9d15476d36d58f1515d48a9ec94a850c121249365d7226fb6aad3a82c9eafe994affffffff58e8d36e4237022b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bd290286ca08485ea4137010c67203c2455e7b669d153c6be40087c7, 232'h0097dd7502ba3637f33baea5b2398647ad24c0fe35072bd963149b5aa0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{346, 1'b1, 512'h792eae16afd3069393b20db2ed2e192ffd845b08e10d076d8eafc98744329d6279d31d55ad56a090712fe131358feb130a94bc4a2fffffffff97daeec1130838, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c917269a5a4ce80b7fe54a8bed49326b50527a4d2fb0a3093182b5a5, 232'h00a195ec0e69e3172e854e87dd651b44433fcd7dcbb7bd59515d2afe8e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{347, 1'b1, 512'h51ae80a63d993770d8a5957111af53dabdf3abb9cf9908bc162ded716d3b3c5af2924c076e87c96249a4d7650253ff5112f8a2e7d2aaffffffff66e0e9175efa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0b7b5aab8364dd4b11001a0b986d5aa4fb61ee720237417a7f63722f, 224'h7f13b411e645e819fed1b925ebe807d9560b44d0ba1b75bd2fbd1294},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{348, 1'b1, 512'h100c883756f36d7c944d934c08932a99a1c2eb9892cc39a13a80b22aadc526ad755265f9ebbc8d0c1ccd31240299c71604332ff56592b7fffffffff1224308a3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h505b974f8ecf07b60ffdbd2b2df9324de92b39476eb763a4c25f126a, 224'h1c36ed1dee772c724205f717c383f49a87a5bc3caa0ef81360f9d800},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{349, 1'b1, 512'hf4272253af2b51df321249280f3f3e62fb1e4a4a556f88bf3d5ae20ac5cc3e035e7b2141f9139b2f21d431068b8d5d96fcaad0f106289298ffffffff51777f01, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h24219e49b98a9b64e56d21c908c870eb88b447d9f1ddb735083d6df2, 232'h00bc4d7644faeff1e134443b2bb3bb2a20e2a4a7c193180626127ce937},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{350, 1'b1, 512'h8bfa5531067a5cbc9bf002be2397bd10dd183d7ae47a02c0d0a7d87e1f94af93ea7365b711cfa611750ac963de0551c900dbad9cd8071b503afffffffffe6b6f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h083246081cf2f8c5e1cd42b60450fc6cac3b0ab03d38bdd271cd7370, 232'h008d117ec32dbf939394499f7dbc2ab77290e9222d6d60ea02ce45c58a},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{351, 1'b1, 512'h8a5409853b325b917b8a2aa1eb394767bb07fa82af11357e777f7404e0955bc9bb9cc5a918475c52df4772a1207e3ee4f3e3d3c8e68e84e10477ffffffffd35f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h24916961dd0d168c2878ca4fd065b81311c03b7f23f8416f4a23b14b, 224'h1e37e3c03b2333b33bbb2ebe05b031042af19315adfdccdfc8d078ee},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{352, 1'b1, 512'h8e38a571ec826b9af00de0c523b6e073aaf9380cc64fbc86755f33f065361d8963ea2c42796ac7516f53d689e1da364bb7caf6b22a5fee81410646ffffffff7f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008df5468b123b92477a5c57ea86c54c5c9e41d119370dc18922aa8303, 232'h0086bdf06b75f4d49d02c5806926f5d01b1a4f6a8146664a03fa820772},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{353, 1'b1, 512'h0f3ad12803aaf9bc615745a47da85dd90bff191d3e9441cc2cc96bf8c01f5e514b256685e3e48f01a98a5f27d20cd1c317a6f816ca8611fbc8891236ffffffff, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f65bf16f7ced97b0cdc22b08c62ef811306813134b001bc51140e828, 224'h3a9b7c008cdaf803368df9ee50e274c7a9f9369344d9918e0c08dba9},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{354, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6239877430e268f1a3ada2c90357247c6ca6687f49023bed0fb5b597, 224'h355c60c09f0dacb9d74b7ccde71806c50fda8750c6ecb7abba910ac7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{355, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h4408e5c95e332ab6c2823a63959391d60a6d69c59eb1f7bd272206b9, 232'h00f5278e901fb4773aeeb2d8255ba4df3cf3db7e0557dbc6134c55f3a6, 120'h00e95c1f470fc1ec22d6baa3a3d5c1, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=120b(15B), s=232b(29B)
  '{356, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h4408e5c95e332ab6c2823a63959391d60a6d69c59eb1f7bd272206b9, 232'h00f5278e901fb4773aeeb2d8255ba4df3cf3db7e0557dbc6134c55f3a6, 232'h00fffffffffffffffffffffffffffffffefffffffffffffffffffffffe, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{357, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h315a83008dba00b351c3f9fca0811c3ae1884fa9a2a75e6d5e71f269, 224'h504bbe6a25be253b582efab4b8b9e61372767a7a3a423c0943127296, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3b},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{358, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h2f6983b6e9f8ef96c2d981f69be54b06591ed73fe40c8a546b936a79, 224'h71bf57726c26c811d7625a9d851951c1fffe236b0eb3b896bc4c98ef, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{359, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00d1f515971cc9391153569c2befa1f915e2931110757760ebd7e61f86, 224'h41c3db8beea20b13205389dcc4ba8a6af4d6da2604cacd7184ec9dbc, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 232'h00bf19ab4d3ebf5a1a49d765909308daa88c2b7be3969db552ea30562b},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{360, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e8f90a717714f0158d9521f18c14ae8c83bf1eeba115c46cbdabb20b, 224'h66f50ac13461c02da02edfe4296a1f543dde7b4359f905e04193d3cf, 8'h03, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{361, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h723bc0c9b7ce6ea784ec075036cede90452c76576bd8fb5be4dc0fb1, 232'h00cf405820d92f48552b551c7b11f49406dc892fd659971ae7f9e74b59, 8'h03, 8'h03},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{362, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00a0dcce127084f955a4e49a7c86b9b91b05ae7afd6eb07225a6541d88, 232'h00f10a1d4fef93934967bb6c5d8792bbd47ab3abb406899a00b1c91b4a, 8'h03, 8'h04},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{363, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00a0dcce127084f955a4e49a7c86b9b91b05ae7afd6eb07225a6541d88, 232'h00f10a1d4fef93934967bb6c5d8792bbd47ab3abb406899a00b1c91b4a, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a40, 8'h04},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{364, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e10abc9fe15bcc63f009e161aaee26602415bcb45bc6c99ce7ab2b10, 232'h00fbebff4e4de0dfaaf04594dd603cee80b5d9ab78b6707608a95e574d, 8'h03, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c6f00c4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{365, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00fbfabe6c640856ae5dcdc9e4b706fb3db23ddca46b80b9057ab9e44f, 224'h6b62d4697977ffe19bf3185083b1ede2161aa5725401a8f57851fc82, 16'h0100, 232'h00c993264c993264c993264c99326411d2e55b3214a8d67528812a55ab},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{366, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h0091a85b3c5e90b409f6b8d3bca9117a54a40f4162b388bb9367fd6439, 232'h00f1cedf20ab52eb7154b7ea1f2934a9c8292906e18a0e572002cd2f7c, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=56b(7B), s=224b(28B)
  '{367, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00d1ca7a5c1aa086b2951c1ac14e005f0072fb28383973a05117f9652c, 232'h00ce523c05ebe94991c47fecd241d0a07e86c88ab3c620eae792aba3d1, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{368, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h3565af2a481f9390e71d7642717d0427e02e5e7de8a3c0c1ffd5f33e, 232'h009474547e0d54dcaae85494c74faa23394a056e41c2839638b8523b72, 16'h0100, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=16b(2B), s=232b(29B)
  '{369, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h29c694790fbd23777cfde434badcb061a326a5534264bcfe193c716c, 224'h178a943f7bd4fb132565ba602358b13433a5217ac04cc035566c73f8, 104'h062522bbd3ecbe7c39e93e7c24, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=104b(13B), s=232b(29B)
  '{370, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h008fd43aac8556f4665fd4c13f4e151140f42a395763c5da247a398f97, 232'h009687d24a9fcd6b20a59451c348a6364d0ffaf0ecfe164313db6594ab, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c29bd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{371, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c2ae0e357a43f97549a725ae3704449051c96bf3633355c35b6eb7e9, 224'h6a84dfb6d4517d1de46b18786a506178724bf4ae4f9e418c75ab17ef, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{372, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c2ae0e357a43f97549a725ae3704449051c96bf3633355c35b6eb7e9, 224'h6a84dfb6d4517d1de46b18786a506178724bf4ae4f9e418c75ab17ef, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{373, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00961617d9855f202fd600b584abe94a46674927cfdc6333c5be56ce7b, 232'h0089b4150d9ccdfbd77e7682ca862c0c3e96d89c918b7d3b7bbb92ff43, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{374, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h008db53fe4168df43ee538bc9d758b8c26fa433fb0101bcbad039585de, 224'h2310dfc20835379ea406993036fd4bb0f67d14760e1eb414c32dd1f3, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{375, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h0b7fa61983e7a227f738847d457f3e8cf0a4085c312fb6dcec822570, 232'h00ee7434ce2ff3fbcc1d0960379876e9dd5bed28aad576eea233a44b0d, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{376, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h55b212919cd6886b13cd7a2556430ce442e86942f1bf6e4618ae363e, 224'h795c664ae960ee1106308b7dba91240ab0c3ef8beb7d0a4d7a102a7f, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b0},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{377, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c0288a63ce32263f3651198dab801c896fb9308362fc40e35959e140, 224'h10d00bd1c228cfb6a5faa647387804e34fa1a7f9fcc472c05ea2eeda, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00bc07ff041506dc73a75086a4325211e696eb6b31da8ff5c2c728d38d},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{378, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h0c8e2cb5f6a903e1cccf3ac2d465f1d0dc3452237fd9e8a4df5d5341, 232'h00d044ca8ceecb54a1b951270971e5ab4eb226116c48c553499d1a4899, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{379, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h1ff6b9901784d88b25527b3702622a2734b83d8a0fed0f740bb784e2, 224'h0e83ee0aa82933dcdc637a3760606a04974c2dc75f12095f8fdaf003, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaa0f17407b4ad40d3e1b8392e81c29},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{380, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b21faca17b68058752d943a81f853b800562df8b2172e150953c6242, 224'h01c2c0f5ed3b342956cacd26f9097562d0fb0a3ddab91c5ae7e90c01, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00c152aafea3a8612ec83a7dc9448e6600ae6a772d75ad2caf19f9390e},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{381, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00f49278419e4f506889b0168b1fce1f87ee5b61efa0e73c7833eeb29c, 232'h00b1b334f81be8f05f3b2e98d38b030cff57947b96135ec4465c5e53f3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h4e158ef86cc53054f1635c74e65508206048929315e097a59f1519e2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{382, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h75c6a886e22bc04b996d4a19575ce0c6686b449b6e05ef1301bd8ba2, 224'h33ab29f65df2d4144da2b21e90359a064765c95e325bb7e54ca28e40, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00e2ac0b24512e84f6fb015620d689d30d14736cf00c18838753c3814f},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{383, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00f554014cc14f319c18f5fa6cd739249075ff35ba3b2afdab5329ef0f, 232'h00d2c501f25a704addbd85c0e022748956e5998d99c387fbfd343c89e0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c5221f3c2de0c6fbc07ff04150679b57f57512b814f413aebafe731},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{384, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00bcfa8db704aca56feb23bd4b4049213233aa652045a0a81a2e0da64c, 224'h091b359f7be7ae00a0e9777d9510f847430b5dfda878e66d4fb0d62f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h221f3c2de0c6fbc07ff041506dc71b5a312063d87beb4c30c289210f},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{385, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h009fd4d828ae98056be58fa69eaf9cde98ca0ed9b415d6463fa1864d9f, 232'h00b2a5e41f10e8789450217daafd259f204aed87b0e26100f43f7c5bad, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h443e785bc18df780ffe082a0db8e36b46240c7b0f7d698618512421e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{386, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h6123a33969f2e036fc27885f55755d391cb0c2d3fafb0c4056c1995d, 232'h00a03bb490047e88fe7e608912a6205b65f950a8a0a360362d3339e62c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00c2de0c6fbc07ff041506dc73a74fd50136878b7e1341521b2f880b19},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{387, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00a10b7aa7785b2f2791b1d4c43e127aab5669612d740b38abaa0d306e, 232'h00c178f216fad379ad80baa0eac57bf9a56d446d685576371b74762382, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h009f56aa80ae2bcf689be2c11b5db7e3a28983b4a7590692edcf5f8db6},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{388, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e012c23c6867e9553313d0179e9db953de7c368cdb59abe05f1c52ba, 232'h00d352a57bb59c45159352c114eeb696ec3b79caa835ef5c2ae71ddcfa, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3ead55015c579ed137c58236bb70b0a2324e79109e2ffc964262f12f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{389, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b9ccd7f0f3594954aa729bda4be883e107e7f1226465b64c2ca71057, 232'h0089829d787016c5c118d3ba3317a2da0a0daaf56d3004c10962333a9f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00de03ff820a836e39d3a8435219289444bbd22db7f7368f8411c27ee5},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{390, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h321a17de024fe89c1864e128b9e0af3e6b48800a70d6e802b8b6dffe, 232'h00b1a8ae96911ddbdeb83948a992b1b0fe316679c64814b6a45ec56fe9, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00f15605922897427b7d80ab106b4474d7fa962e970ffad666580fd5c6},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{391, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h08842f19b114d16be27bb4b6971377ed6b1d0915e133a9ebf01674ee, 224'h4c97738b6912ff71553c4a747c782eddd9d2a20fbeae38864d217859, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{392, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h0084d651596fd2348f1bb5c8ae9d22c8b21c4f7509240b609abad5cc24, 224'h3196b67b4cfaffaf0dce25ab00bfeaa1a64821332efa6dedd87cc9e7, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00855f5b2dc8e46ec428a593f73219cf65dae793e8346e30cc3701309c},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{393, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h008fbe39e75bc4fd8a15e4b52e4bbebe2047d54385a7117e17a4d0b2b2, 224'h07abdb40824538e5787c718d6548583f523f6b5bbfa239a7f622c8a0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{394, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c336b340bc99d46c2c52df5428b6a0c4eb2da76c423530f767cc7652, 232'h00f3ab9981bd05d2955123935a379cbb2d4361a17d19878673e1e17dcc, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0084a6c7513e5f48c07fffffffffff8713f3cba1293e4f3e95597fe6bd},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{395, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00816fdcf370827e3f7771564e1aa73ed73e62556deadad89711cef663, 232'h00edcda0ea42235f4c9a8c13f787351ffe5ceb32f15fc0ccb24e0a409c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{396, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h6429d2b7b07ab0d5ea352902df0efc036d7270a0a6ed39f635d04f39, 224'h4f7932883bc45394151324aab26ae29bbd7385fa6a42c3db84432897, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d8ea27cbe9180fffffffffffffff3a43fa3662a899627950d4eb64bc},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{397, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h288f38fd77dd1603ff0275cb11cba280ae3408affa6a760f396f1a1e, 232'h00c84ca6fd772c6ac6cc523cc72c2e7e95eb6a36a66b5cca5a58ba078a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{398, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c769c138f9d71ffff113273b71a4afde4f9996a1c4be658a3903cf7f, 224'h430e512b868b37bb96bc17a09b0ab01b262f2e23f34f00418f6b63d6, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00bfffffffffffffffffffffffffff3d87bb44c833bb384d0f224ccdde},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{399, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h75f007c11b93e6f46e9a815cb765990a8305d3ad8d22c76fe6b257cc, 224'h71b5c1951b5d464c66df7c290cf0a4f156bbf52f1e41a79dc63abce5, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{400, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h1255fb94a0f20e6faa2505c394cc3c39f07def4107127dffc4dacb6e, 232'h00ea73c1044544a1496560bd1b049ff615e68ae0d483220327569884e1, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{401, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00f656a632a0804cf688446b261208f793373c5ff4454bd1e0a882113f, 224'h30a25d6f586e02dd4dcbf73d96af3e483b7acb5f8f4c06450dec1982, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0096dafb0d7540b93b5790327082635cd8895e1e799d5d19f92b594056},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{402, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h008fb572de4daf76702624ce4ed819d026762224e8a54215bf81b202a3, 232'h00f074d20e1da7232d279461732bc1bae0c5416ab9d696308622e7ffe8, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 232'h00ec0ce3fa725c1027475a5f5bf4ee980de61c3b4875afe8b654b24ee2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{403, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h008fb572de4daf76702624ce4ed819d026762224e8a54215bf81b202a3, 224'h0f8b2df1e258dcd2d86b9e8cd43e451e3abe95462969cf79dd180019, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 232'h00ec0ce3fa725c1027475a5f5bf4ee980de61c3b4875afe8b654b24ee2},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{404, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e5462d3a838d4a14de96a7b0b1071eb622ae6e71ede8f95ff01c2121, 224'h368e3a90d8584e194616d3211a7541f6a0960339cab28e8bfd6b1dfd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{405, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h5d97670c1f121f7f1ba541505609f20143b312a7bb49d376690e1831, 232'h00c1b4567141a7b534e21bd2f706ae034169ab9c3f8536147904de8c5f, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{406, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00d2675278da2d7daa8373dd63b7aa46cb14766571c2d8098b83a102a5, 224'h699b572d4b951497418a376930022d48fe59966b158fa08340e24b98, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{407, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h5a5cd1162388348734dae20e2235ae2c464adef0a196f9aaf02482ca, 224'h2ae94e8b9a024375036429b632ab485e02c5a9665b289b8a47bade8f, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{408, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00cacd93eb11a821de3d882bab7411e7c77f23c08da174189cc987dc41, 224'h716fe378ab842161bc16def6e037d4ba9d30d8cb41ad30cf0656e50b, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{409, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00cf46960060453e55577f1bee6a9c4709e7cdcba45ca8020bb3536931, 232'h00ea4ec33309213864a1318aee0a86d8b6f0c1b9741cd6bd5dea4f4066, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{410, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h62f4eaf3797bdc3d5d8cfaa07b5af7060e131b183ca4eded4819e561, 232'h00bff3eadd7b55db2dc01bd20569e6c47c9212f9b2d6793795b51e4f6c, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{411, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00c4a4bf5ae0138587f50ab7a2c336a430527a86f59f9765c2f3f5488d, 232'h00f9419bf9df5f121de3a32db17b49c72b606b2be5ce56acb565cc12b7, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{412, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00e7cb5ae54dbe619ab5069f14566236b3c6b0b44f1c4c531e66d89b3e, 224'h64be7fdc18789629dfddf7158f8ff27abd553bfac3f7c874bccdc31b, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{413, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h30db5d8279319cf5a3b6768a0c5e5c84752f6314f735d63f6c5650cd, 232'h00d32fb54f74d4a5088e6774a13201683642790d2e69e55e4f47612934, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{414, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h7db27da4d67a2de0c78815809719bdf6976332c67ef0f3827df4adc2, 224'h2ab37aec2eed0d5e67acfd6a195f21032d9af71ce73e120fdda29f1a, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{415, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00d1c19d46b517bb3bd7bdf074ff975c0dbd2bde10d1ad217e58ebc8c5, 224'h5ac898c040a185804ddb032b48103d6c8d12043d3a4fec93aba7a6d7, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{416, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00d95ac96ae9dbfb80911862e00a4cadbcb2359f499b53be007f0711c0, 232'h0093d3da931acbb9242800dc521695b4f19ff2dffc3613f40bdb15c3cd, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{417, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b0, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{418, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 232'h00bc07ff041506dc73a75086a4325211e696eb6b31da8ff5c2c728d38d, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{419, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b0, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{420, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 232'h00bc07ff041506dc73a75086a4325211e696eb6b31da8ff5c2c728d38d, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{421, 1'b1, 512'hcf83e1357eefb8bdf1542850d66d8007d620e4050b5715dc83f4a921d36ce9ce47d0d13c5d85f2b0ff8318d2877eec2f63b931bd47417a81a538327af927da3e, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00f72915d6d916014279616186869a01228fcd9f1b4078353018b399ab, 232'h00b67f2b91eeeb910381f5b461a4a39c642aea4792013d4eb63da1832b},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{422, 1'b1, 512'hdc5e71048a56da7aa1bf5fad1ae227446663488d8a531d490c4b5efa048ca4651acd9a196d9b13ee2a1c74ad440bdd88f6a34a02fbfadac2f7ce869e64486558, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00a5d179c336ccdc760dfddd913cdf8ea468d0f4686f7b2d3825698ed7, 232'h00a77f12060a4d1b94b0d1c443eae3ad6e21b7eacfdf6fbf39a2b29658},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{423, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00b7c65dce56abe24fb4592ece5ac1e6ee8353431f7452409add736884, 232'h00e5fe5db7988931026b937dc4ef983fe446ca134d29b94ac777cde317},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{424, 1'b1, 512'hd296b892b3a7964bd0cc882fc7c0be948b6bbd8eb1eff8c13942fcaabf1f38772dd56ba4d8ecd0b626ff5cef1cd045a1b0a76910396f3c7430b215a85950e9c3, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h05c563d3a4bad874e4610adfa57777a59f995bfa06ef97bf125a4988, 232'h0097ed68f546cf4bb4998524c18356f3af162d2bf2744be93357bc4b4b},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{425, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h00c7a6f358b7d93815189ae5d2c3ab4d4e05f43176a52dd4fc5b48a34a, 232'h00a2458512bb8dbe6f1bd6eb01d2d77d5624e8547bf87d85fc731c0c86},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{426, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h5f56ca587d16664a20dad13df85a475978e5cee81a8d0f49faaf6158, 232'h00b64ef59d79461fe1a09a5864907435f70bd75f183afb11903f560b7c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{427, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h00dd94f5b56e9947d007e7c8efd894a5c882f1d0b5dd56c32b5b266521, 232'h00fbc883741bd27c59958ae17ba6e4a41ad1edeca9a3ba31c8f233b5ac},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{428, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h008071e6682c6e8a32706dc7e411503946546b31fff27dcce188ae389f, 232'h00dc396c797d44edf794432d1da091f8c762974d8ce1f06e08ca013622},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{429, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h791624e5f234b8950d509d0b456ef6fa778b19dccd609d496b62a211, 224'h6c51e846fa53d03d42f798e6bb90954f9a48c1794b47e84ac97b460a},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{430, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 216'h34befa1d25b756ce76b383a6e8753741c12a59266c2c7921ff6e8b, 232'h00bc44e3823e4d807cbc92fa786a89e62a4b217b5fb0c0f1865d4a7e43},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=216b(27B), s=232b(29B)
  '{431, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h224a38e733ebd3fac274ecc50ecef2e7c3189be2b9d093a8dcc6fa3a, 224'h134fa5a4f923d296b3c6dd4683d249ccf0ad272890e4149c9a0d7415},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{432, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h338d07d990879ad844e24c1788e362269d8aca70500357d385768227, 232'h00f745cc4ebaaf1cd42830026a66e5b95564cdbee5edf853bb2cc91259},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{433, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h689fce4b33d8212a663640a1ae0efaa7a7d7711beba719374fe634ee, 224'h04bd9981fa52293063076f0fd70fc31875d580ef94f020d2f95440e0},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{434, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h2a4287e01510e7fb5fed2e1ccc3f2a6929cf7d03850e49d7ae8a504a, 224'h355c3915f3fa9637dc8001438a8c04e15d14934cabd430feb0cb5ba5},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{435, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 232'h00b5bf795a38adb052b401468ffcab81103d2d9fca2e15b8d08ab98ce8, 224'h5ec0d2c6aec71888c941af324c7272bec192abb292f9df82a24e8a41},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{436, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h100ed07f467133bf10917f7a15ab2bfda519bdbc2653b95955e22211, 232'h00b38a081f7c2e2b775d1da868d0381c09ba1559c9613b5be7159363ad},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{437, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h54e6add8ac910e52c6228fe3980d8f586218334d8d859ba9a3329917, 224'h5836cc79ec88519eab4a6b2614c501628c9fee32fbafd93e32158409},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{438, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h1230d5409f379584b4d548b7bccba64baf81d512a9f2e6398c4e3a66, 224'h1937a298f8cbdfa85b8e6fcf0a12be4966d80270cade85a0c37ee6f3},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{439, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00862f43b044fb32adb45e00378ba083ae761c84452054f17b1341bf5b, 232'h0095d8d8e5e3a6cc2b0a06c792252ca11a642257721831578520f96b9e},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{440, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 232'h00cb5cabb1ca01b847a6bc70558d1e5d3a204d1741bbe800f4b159af35, 224'h3580cc85f218394130bddf1c4eac04fe96f59f14fb436686950398be},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{441, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 232'h00c9d83dc04cf4ee89c405045d0fd1d704f627ca5bbe350f40b826bbc1, 224'h74fedc9e55045e9759f2124460fdfb991dc620cfee6effc0b4adaa9e},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{442, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h46dd65b6e7f10c0841841b01033a5befd3a0e78c85f1f390bb3cdf25, 232'h00f33acea3d47cf0dd5273735b004104f6512ed641052509422c0325a7},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{443, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00ddb4a7e400a1e98118f474722da3f421f65a76eec61f4f7b699faf07, 232'h00db80cba199859cdfe916d6ab3deb91d76aaf0ed554c8f9ed7e5aa59d},  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{444, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h4c260b546280604e4c80384721c9e803ef704e7fb70168e6730fc1f3, 232'h00a8aceae219ac25c9f04231b4e0c171413db1d26df1c1e8430062eb2b},  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{445, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00f4098d2c0240e78fceabb0183df0b39e7ad3e7f5d6da1587fa09853c, 232'h00d42412b2abaa614c95eb11f9b9346282ce3a1c93aac35ce7aa372f4a},  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{446, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h48ddc497f9a4732c677e46c0e2bdabec54fc9d27e46ab595056db4d9, 232'h00b8219ebbfaebc2fe4311efab0c35d4392751351bcc1971e8d01941e4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{447, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00e1abaf51d27a6d7d4c9b28078325cac2d7ce3d5403916c68903760b7, 224'h2c45a99e2770f782fee5ca1d713eaecf07e62d53c64b7cf93de9900d},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{448, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00868cd127c99e1149f7fc8d878cdfa986b62e99addea281149611ff15, 224'h16e5953820135b7d462ce5434ef85920e973eec9e4d14d7cb3cc2a3f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{449, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00a375929718ec4e6ada9c9370c51df6bdaee7ebab2a70675d42a0b6b3, 232'h009eaf4802efaf7ca082ffbf5ed774af43792d9b3fd711c6b1c36112ff},  // lens: hash=512b(64B), x=232b(29B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{450, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h00d97b32f3bf8bc11ec2672dd6320418beeed99527a63fe4c52199ec61, 224'h68dd9006b03319ccbe651d0bdaf84c63356f03cb007a6865ee3e0206},  // lens: hash=512b(64B), x=232b(29B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{451, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 232'h008ee5794dc2e66f2584910ea1d8361e5b53db535adcf5c1c35e128309, 224'h5d1d8b9b996c0a488e05af14421b86e9841f0cba706027fc827d4d95},  // lens: hash=512b(64B), x=232b(29B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{452, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h7999727c0cc02d88ef274012a762afcbb19e7fce19091a02acd00564, 232'h00dbfacf67999f22c499d48a60a6fe4bbb746199c29957a1ec7a0900e0},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{453, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h5797c21c0162e42f69693c6c0244dfdf9218c01e9235760177b61a54, 224'h5452c887b27fb342a8a00d27579c7195dddb73df399233ed0dea567b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{454, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h0eb9dc5d67bb0d4009544f8654977907dfe770e7fae4571d31d7b4fa, 232'h00ab5cda53e868bff5198be4be3681b186cb0c1396d272c71f093f8b12}  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
};
`endif
