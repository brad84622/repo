`ifndef WYCHERPROOF_SECP160R1_SHA256_SV
`define WYCHERPROOF_SECP160R1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp160r1_sha256;

localparam int TEST_VECTORS_SECP160R1_SHA256_NUM = 230;

ecdsa_vector_secp160r1_sha256 test_vectors_secp160r1_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'h00a064880a1352852176abfa15c2787c05d84f5e8d},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'hc0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{3, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{96, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 184'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e50000, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=184b(23B), s=160b(20B)
  '{97, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 176'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca0000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=176b(22B)
  '{101, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 184'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e50500, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=184b(23B), s=160b(20B)
  '{102, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 176'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca0500},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=176b(22B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 0, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=0b(0B), s=160b(20B)
  '{118, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 0},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=0b(0B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h02c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5d9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff2965, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c34a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 152'h5f9b77f5ecad7ade8955fab336af32cdf225c3},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=152b(19B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 152'h9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=152b(19B)
  '{128, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 32944'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e50000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32944b(4118B), s=160b(20B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 176'hff00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=176b(22B), s=160b(20B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'hff5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 32936'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=32936b(4117B)
  '{136, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h01c0d64c9119a1ef31b0b49ad41dd0e4547d744c3c, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'hc0d64c9119a1ef31b0b0b1422b8186ace88a078e, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{138, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'hff3f29b36ee65e10ce4f4d59f4db56ca7f4d00d61b, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h3f29b36ee65e10ce4f4f4ebdd47e79531775f872, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{140, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'hfe3f29b36ee65e10ce4f4b652be22f1bab828bb3c4, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{141, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'hfec0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{142, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h013f29b36ee65e10ce4f4d59f4db56ca7f4d00d61b, 160'h5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{143, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'h015f9b77f5ecad7ade8957ef7c2fd6e1a1bc9ae621},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'hff5f9b77f5ecad7ade895405ea3d8783fa27b0a173},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 160'ha064880a1352852176aa054cc950cd320dda3c36},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'hfea064880a1352852176a81083d0291e5e436519df},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'h025f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'hfe5f9b77f5ecad7ade8955fab336af32cdf225c3ca},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00c0d64c9119a1ef31b0b2a60b24a93580b2ff29e5, 168'h01a064880a1352852176aa054cc950cd320dda3c36},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{153, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{157, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h00, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{163, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{167, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'h01, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{176, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{177, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 8'hff, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{180, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{182, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{183, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{184, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{187, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752257, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{190, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{192, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{193, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{194, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{195, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{196, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{197, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752256, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{200, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{201, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{202, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{203, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{204, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{205, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{206, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{207, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0100000000000000000001f4c8f927aed3ca752258, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{210, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{211, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{212, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{213, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{214, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{215, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{216, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{217, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff7fffffff, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{220, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{221, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{222, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 8'hff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{223, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 168'h0100000000000000000001f4c8f927aed3ca752257},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{224, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 168'h0100000000000000000001f4c8f927aed3ca752256},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{225, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 168'h0100000000000000000001f4c8f927aed3ca752258},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{226, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 168'h00ffffffffffffffffffffffffffffffff7fffffff},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{227, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ffffffffffffffffffffffffffffffff80000000, 168'h00ffffffffffffffffffffffffffffffff80000000},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{239, 1'b1, 256'h35b67cfb1515c415dec6671a2010bf1ef24faa0518e5ec635aa7e3cd0640c53c, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00de3a6ee112b425f2144e452abaa9d11a237cec61, 168'h009c406f41e1688cd89e0a1651c5740c961c59949e},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{240, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ad3f5fc09120df90e8740111934bdc50723172a1, 160'h410ae1236da5eda0b327bdbc9e6d545a34764051},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{241, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h2a08a7f52a3506c5ff0b0bdfc41ed256a998deca, 160'h3d5324b851f80f334befa39b77241cf06535a1f6},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{242, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h48dbbef868af35b058bd34e507e85fc61fd60f31, 160'h2efb7e448ba59de5835198c3d5f5015113a3dae5},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{243, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00a679ae2d7bc1f7d4c03fb2325928b253b090a56f, 160'h646f90a9210a87b28324d7c50a454abcdca7f53c},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{244, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h47398e906863d57ea273977083d36ce35f1f619e, 160'h24959c9b1f06bb8822bd8fac8f45945fd1c7ebeb},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{245, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h599bcba0ff3fe6f2d8b2544e3b824731666d19b1, 168'h00f5d15469fce1e244750792f327bb6ee5e8299f94},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{246, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h4b24155af66bc983050381c2579ad91a85c48d4f, 160'h28b0d445e93fa372a59b7030c67d2124b9bbd65f},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{247, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h57999b6dcf7d77337d8445543f1ee0d212d7f85b, 160'h5f4c8fa2f113b3637504b42160ddae852daa1d78},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{248, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h0788eca735904e004f414f5bdb087365fae662d3, 168'h0099e52af8c7f20ce34f31831ea32f6503c03c3a29},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{249, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00f7bd7de59fe7791add20a4992425e20c1435de4a, 168'h00c5a9fea1317a237486a19894c4e2e8475eeac5c5},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{250, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6e3647dfed9c5ae3cc481528a35f5741e9dc10c1, 160'h569c3937c0a118cb49358a640670916ba346db03},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{251, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h5f603ecbac6982960efb6d8853de3ddfb4b2236e, 168'h00b4b779028c7e8ea850242607e6463884620188ac},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{252, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h1da6db19788b81fc3ddb980bdefa9a54d33717d0, 160'h018b151eeb8c79bf5be669f12cb784615e098317},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{253, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h7add46bab0d2c221d03f6a93d0fcc9e1a54b0c72, 168'h00b1781bd689a5334597b802713a0fd6f561132c82},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{254, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h008311662f6c665414a4eba51c328b0379455230ce, 168'h00bed6cbdce059464888cb4912aa34b5dcb9e62123},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{255, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00f86aa3566274a62777e474e85598fa2d56ae19e4, 160'h459c11cbc8a2ed4b794b6deed3c7ef7a4a45961f},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{256, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h3c2c6830a0733d25facdf0048a9d6c3b2921aecf, 160'h0c7e0c333dc82930f5f8a4337b379db7f0a526ee},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{257, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00face1b45e18a0f9dabed5ff09bb800ec0536987c, 168'h009e60b1c0a87937fc198034b4365622290cab54c1},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{258, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00e3cafaa1fefe07ba010efe4ef7823cbb2e05d32b, 160'h151f1b481a24ddd5df98c04d058548fd06f47f21},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{259, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h009bda6733d547555fd2aa1391ff421302005d2a4d, 160'h4aac3e7c1dbc99a85560a921f34ecb3e8ba37466},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{260, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h53a8f7b311fbd2b71cfbc781c50923bf4c423335, 160'h33cf2cf617f565b831d82e93e8fb58de938dbbb5},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{261, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h3332e2dd4080616b964e7bfd569e7b3ca0767b38, 160'h65e0c755d4dcf460fbbd2640d347298f2a29c156},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{262, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00d94703055d7a99e1727c20182565339945693cee, 160'h0130502398839f604729760999ed64350e576517},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{263, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h5c1a34fcc2cbcaf2778e85e94ada69e18ab40648, 168'h00c3798cb473af1d33b2df5ddfd7d48329dba04d31},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{264, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00e063a77c688cb1a3deae3cfc44b9004105aa3c0e, 168'h008f1e9b2fe1239931b0aa35b8ff7d555f076e8eac},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{265, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6f11c31e65689b848136fe044722081ded5f3bbc, 168'h00e975164548bbaff051e8fcbe3e7fd1da7460527a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{266, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h008ec112600f5423fec61a9eac11c2d7f202660afb, 160'h3c3ef6efda5343622a9cb37114989019bcec3016},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{267, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00eaff9d359729732e49327affafe0750e42be994c, 168'h00b4f2ec9b4ab9705c1e407ce062b4220f74cb8209},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{268, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00b7237f113c3c39892e21bc1530089eb2623e1ab5, 160'h1647796cd696dbf9fa852b14ee59b103823940f3},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{269, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h41d8153033a3144823afc2301780de5cc70792fa, 160'h0a9add978d502c71a16a0432451513c7255a4ec4},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{270, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h0094b7bbbb637080eadb0052b09edc4e1cf971af18, 160'h3fbe47451bb32f532c4f7c87125d40bd535f4478},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{271, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00eadd4b4acce3825872573405025d1603eea896e4, 168'h00df0a9702fc9e237d05ba8ffdc37f646df9cbebbf},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{272, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00a5bc403170737f5f296da2edf46c979b00f6b4bb, 168'h008f0ce6d5f7e485753bf3f850254c5c32b385205a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{273, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6f10822c847280ca0c687e209d7738db57315dfc, 160'h7ffbab843768815a87be79b2f1edce6be8423480},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{274, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h40a127c4d89b3e793bc7e42d3931266e2e2b7acf, 168'h00bf18fa3b5982dbdd02d4814f5a0327fed477646b},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{275, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00acfc8f05a71e19aedd5619453c827caec3e08204, 160'h4163d41bd88c689114bebdb0b14ca63de2e636ae},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{276, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00b381bbb8746403e6fe9d77791bf6b9ad01b8c32b, 168'h00e793bf926db9c1ee35daf0457e890d34e3f702ec},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{277, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ff086f8fb05d39d6718bc58ad004bdb1a3460e8f, 160'h3661b0d1b65b20f5a6e77aac3930b08f99efccd3},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{278, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h009a6ac4de9b691f5d8e7b8620e432672014dc14fb, 160'h19ed53655eb2795b2e44c1a69be207e5a12f94c8},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{279, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00de41eab8fbe839db07b3aa27580d87fb21b0043d, 168'h008e9b72997d8ab82a4c7391d94dbb4904231539b0},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{280, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h40bcf243c5a448103497a72ce415850d86f9417a, 168'h00bec384be063e3a32be528abb64f8754c5934ad1a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{281, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h2b81c2a07a21637df18094dae7236476211fa251, 168'h00e94a910c43c29f347cfe87cd8cec7d924abb8582},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{282, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00f41ce5f7d5f448dd918485bea20a4a2b7bdb894c, 160'h0bb4afabf1af4bef661dca6573f4cbed564d5b71},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{283, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00ee1309c51d9bb6dff0fd6e182dc910e90745651e, 168'h00b06de7056a70a8b41efa496c4ed4448a423dac20},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{284, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00d74a14b7d315bf1ae536d9f28861eb34f16c6691, 168'h00e7cafdee9e360da3b139fa6b1855391bd4072dbf},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{285, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6b7b7ebfcc4acfcb41a8a6a072b745f274382b76, 160'h38a09a2023d79b6242185529aede41eba8f52332},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{286, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h7caa1b32fb6a67b204878b3694699237eccd0558, 168'h00b1701539856d9713d3eafb326ca181057c781f60},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{287, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h7bf85d33ccb2308d51017419197e53f24a482f6c, 160'h591cbb3ebb4f1bf6571f17b86d07e5f80c6118e9},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{288, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00f876e72b8bd7b156e7ed218186a355a9240c9451, 168'h00ab7df020cbfbf2b8f267290efdf39bc9014558ce},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{289, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h009f6ba902a1ae32d7fb6c62f84013365ca6f9b712, 160'h4c27061486ee0e3da5da9706d8927c37eec8f057},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{290, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h2ad7961a2515241e9d8675c05aa6fa1488714a38, 160'h17dea0a256ab4e20c9554c5f5b0c491271fb0689},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{291, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 160'h6dbf66690812e4bf295181b1c5ce381e9979e6b6, 168'h0080eb3c881c7c8452fe722b78ec4e0d3788c476e7},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{292, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00e2386217f55b3b7f7710d487cefe7940542737de, 168'h0090367b1ec7be80868927fde3d1484a80c4f1a983},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{293, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h009562a2ba7e709d09c6d5daab76a27e14978dc9d2, 160'h15e896d5ce8c1b1512eb033ff1c008d04b4b38be},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{294, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50cd6584a80522992ecc20c20280c358c15e5085, 168'h00e0a12cbbb20fbec12ce194c0f90b72331db90fce, 168'h00a2e4471c0ebd7be819fcbe6480583738c7337e1e, 168'h00bad0f1ced7e0d0ab01adc1371c66e9cad153928d},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{295, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h009452cac89fd846036b3f4ddf995da4bc958e1911, 160'h5f8b30d6cca6988ab496ff2f17e24f08faac75b7, 168'h00ffffffffffffffffffffffffffffffff7ffffffc, 168'h0100000000000000000001f4c8f927aed3ca752254},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{296, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b005b80cb0733576bd27520bf7ac44f28e733718, 160'h09738b9aeb21252938e9a5fa885a4bfa3705e084, 88'h01f4c8f927aed44a752255, 88'h01f4c8f927aed44a752254},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=88b(11B), s=88b(11B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00f0a6c8100e5720ab62dc981061abc4add9a1933c, 160'h3673d536905fbe48defe2b2a8637f38f2e1843c4, 32'h7fffffff, 160'h17644e8c2ec89d185d9167f301adcdedae3f5b35},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h711d5c4035baebc8e46bf09434a8aebbb0f678d0, 168'h008f66aea6922e491d02960c4e1baa2c22bcbad408, 32'h7fffffff, 160'h749adb63d26b6d8f49ae9a5725ade8880d9c9b6c},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b3e8857e27393fb609bb7e4d42bb612704d9eef2, 160'h668439313310a849e17faca660f5f5346e11c1a9, 8'h04, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h1b66bc474c8220de08f3db0fdc984b008828ff5d, 168'h00f94509a6596f822f62580acc988bf962ef9e32b8, 8'h04, 8'h03},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h008ac14539432e062ff2b1f6086926bfc87e342e98, 168'h00bdc182b2ec96ac855f1057cd99731a054067a153, 8'h04, 8'h04},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{302, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4a5c77d11ddaa568733d8a6cb79b497e6a644944, 160'h339c2514eda2e275ceffb9a7fc4c8d0470b37638, 8'h04, 8'h05},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4a5c77d11ddaa568733d8a6cb79b497e6a644944, 160'h339c2514eda2e275ceffb9a7fc4c8d0470b37638, 168'h0100000000000000000001f4c8f927aed3ca75225b, 8'h05},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{304, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h44bce6f9cc091008e68a1764c1eaf56f6fde9234, 168'h00f6bf9770268c9dfb0c2ea33819a7936ee8d57333, 8'h04, 168'h0100000000000000000001f4c8f927aed3ca87f8de},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h5094345ff85c68fe99627eede704362af196aecf, 160'h53499a272ceb4668c02b4b11e567eae9709f0618, 16'h0100, 160'h1c3870e1c3870e1c387118f7eb1684277916fdbd},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=16b(2B), s=160b(20B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h5e2bb1e908df355fb09ac567021edbc0d0fd7047, 160'h65ee7405ef872af6f2550c123826058ebc8309fb, 56'h2d9b4d347952cd, 160'h1164a61fc3dfa342ba186e32381b34b324117a46},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=56b(7B), s=160b(20B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00de53fcbfc744edfc6be04af83518829b5fa63016, 168'h009fed2940a16623e8f60eec87c32aed905d25feb7, 104'h1033e67e37b32b445580bf4efb, 160'h4cb34cb34cb34cb34cb3e2bdb53bb3e1d213282c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=104b(13B), s=160b(20B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h366bb0c1db172c0da7a94d6b962b2bfb99db430d, 168'h00adb55cacb92dcf86d7e7373db40159c23c6ad8db, 16'h0100, 160'h382efed3dc7e18cf41aec7248f4e56087f9734a0},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=16b(2B), s=160b(20B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0086e01061fc02e52057346370636a5b5cc3710e72, 168'h00ccfb1063a51118d442d5044cb0ecdade51ab7dd3, 104'h062522bbd3ecbe7c39e93e7c24, 160'h382efed3dc7e18cf41aec7248f4e56087f9734a0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=104b(13B), s=160b(20B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h40e16716c249fb4743fc761afb05dc34cd447fc8, 160'h179c76ae7ac1f0b0c5f248bdb8140b91ebfeaa2a, 88'h01f4c8f927aed44a7521da, 168'h00aaaaaaaaaaaaaaaaaaabf885fb6fc9e286f8c18f},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=88b(11B), s=168b(21B)
  '{311, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h07970e499d36b850864ce1d6b00d62cb70e2d2e0, 168'h00e30d4b3c346017c766878f93fcbba65cd80a1f59, 160'h55555555555555555555fc42fdb7e4f1437c60c8, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h07970e499d36b850864ce1d6b00d62cb70e2d2e0, 168'h00e30d4b3c346017c766878f93fcbba65cd80a1f59, 160'h55555555555555555555fc42fdb7e4f1437c60c8, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=8b(1B)
  '{313, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2b3a7058fdbd423b96168d487e072feb1a0544d6, 168'h00b6b31631ede8673761d6d3e48e8e966479c08fc3, 168'h0080000000000000000000fa647c93d769e53a912b, 160'h55555555555555555555fc42fdb7e4f1437c60c7},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h59611a33fb3425881e31e0f61f2182e4fce3bd89, 168'h00c0291abfc4d1145a5001de56bdfa96be446d30b6, 168'h0080000000000000000000fa647c93d769e53a912b, 168'h0080000000000000000000fa647c93d769e53a912b},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{315, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h31eaca167a3c657869e55d7e48bcc525c26e6277, 168'h00cf3b34543a52b1611717d94ba8237980ab02e218, 168'h0080000000000000000000fa647c93d769e53a912b, 168'h0080000000000000000000fa647c93d769e53a912c},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{316, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h67883840b961f31142fdaa4225d9186894d533ec, 160'h648886fef0e60348e90621f6b7a553f05d8ff5a7, 160'h55555555555555555555fc42fdb7e4f1437c60c5, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2bea5e4da06c9e290a65d59f9c44f0149616d9ec, 160'h4b9a64a3835d7e249f969d2ccb997878efabaa19, 160'h55555555555555555555fc42fdb7e4f1437c60c5, 168'h00894b5a17a0c6db3c257d25a6ca0a19e1947c7528},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b1fc10305d2e83868c9e40e8426896297b7f3e00, 168'h0091a1e1f88d1fb0f95380f19c98f55a0854c6b494, 160'h55555555555555555555fc42fdb7e4f1437c60c5, 160'h55555555555555555555fc42fdb7e4f1437c60c5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h009eabf3380b193e547dd2610152ea76048806b9e1, 160'h413a8a53711c915d17c16df98300ee414f11dbdd, 160'h55555555555555555555fc42fdb7e4f1437c60c5, 168'h00aaaaaaaaaaaaaaaaaaabf885fb6fc9e286f8c192},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2b9e690b79e165b04e0df6fc84e58ac94ac63a92, 160'h7a9532b9ee40bff794f9888b1a2e0b8a30f4f550, 32'h7ffffffd, 160'h7ce6e1f81fbdb6ebf382414e62c1c14200249a82},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h409c92512c25d7fdf331487d4bb1ca8312ea27b4, 168'h00db6909d4a0768e609a52064c266e152a36b49b7a, 32'h7ffffffd, 160'h304d26aa02922e73b2c60f12e7f288b0b43f3783},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h39226e3be69faee8861f1fbaf4523da7bd2d1bcd, 168'h00c7a528956daf7f7e5c21288732c69372ca327ecd, 32'h7ffffffd, 160'h2b9afe309194473695a328cfe89a314ee772f616},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h74a34455bc9222dc9f189672e0c72cb3d7bf8491, 160'h605793269a796edfb97deeb50f30477571c76d32, 32'h7ffffffd, 160'h0b63c499d27b74e8894b705f6dcab0b5834c4785},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b1031e0781fecf813633cb3884e930913e65ba5b, 168'h00cc8860779ca7e174df787d66f671a8fa337994cf, 32'h7ffffffd, 160'h3c499d27b74e8894b5a1effb88d50da2d531e626},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00987ff07d407ee7a41a65a7ac6929c13d0a6e4800, 160'h59813e21d5f2fe748f06be7328a9862af2bc7c57, 32'h7ffffffd, 160'h78933a4f6e9d11296b43dff711aa1b45aa63cc4c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c071a26e5e5257fe26bdb8013f48bbae17a2f319, 160'h2cf253cf4973d3c2dc250ec4c1e71c1ed3653786, 32'h7ffffffd, 168'h00d27b74e8894b5a17a0c876fa832050294d0ede01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=168b(21B)
  '{327, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00db3da2a11095b2aefd141f26c9b20e43a1f4cecd, 168'h00eb2666f06ebfcfcdfa3f9890769b0db3b85a8a3f, 32'h7ffffffd, 168'h00b080eb3eba27e3743ee6c3ba1d023f83c7643e58},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h0f9d71fb48e807f2e66bfdffab87c78d24cf2d65, 168'h008125943f73180928436be5db4228efb72769021e, 32'h7ffffffd, 168'h00eb2eda56a5606183576c3f3be8b20e9e1fc45dec},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00feaa6f5ba970d904fe254dd45cf4f1d397f8b5c6, 168'h00dbcddef5385bb2ec2e5844b4566cc22f015d864b, 32'h7ffffffd, 168'h0083191e07e04249140c7fb37a9665ed91ca5087d5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h52c0322e296d02806a55800e67b9334ed4005cd1, 168'h00f60f5556e7563b756d8a17cd6977cdde16531660, 32'h7ffffffd, 160'h44a5ad0bd0636d9e12be92d365050cf0ca3e3a94},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h50c07170fdea6845c09c3da29cc8ee6700592919, 168'h0099d3cf10ef65514e890c056a08c505ad13dbfe03, 32'h7ffffffd, 160'h15cd7f1848ca239b4ad19467f44d18a773b97b0b},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{332, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h05cc25d16018b88388a41cfe3547ebda232de5eb, 168'h00bf2017c6bc837a738dca9c8e91b3fbe06d154497, 32'h7ffffffd, 168'h00aaaaaaaaaaaaaaaaaaabf885fb6fc9e2b1a36c39},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e2cada2f22ae694fee3a3287ce8dc0691af40c9f, 168'h00f6a592e8c723bec635a76c9c6482d2b60dddb986, 32'h7ffffffd, 160'h5d0e82e246fc758108ac747e6f91ebfc3800d367},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{334, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h267471b41f818bb8176e2a012f963cd9b6fa2575, 168'h00c14ea6247c7431a05fd7422de905afdbc6c8e166, 32'h7ffffffd, 168'h00e6ae9daaf56f8b83815b6de2e022c30a5fa4f229},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{335, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h009ae2a06f674401b28a799181ad23badd115066d1, 160'h3430009efd1271ea1962d35effebfdf5c94d46d2, 32'h7ffffffd, 160'h44bdeb62114743cb00008678e702d02fe3b75eb7},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d086921c342ee56be74e87950e1c260b070c7469, 160'h0c5ad644b7806b75469af63d8ba276c568e8e27a, 32'h7ffffffd, 168'h00deb62114743cb0000001b3aa8fa7770551110483},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=168b(21B)
  '{337, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c5f85f1245c93cf37f8258d3f18e15ae64bf3724, 168'h00c3c3f7dc1229fb8b5ad0274eae7c98d5fc9ef67a, 32'h7ffffffd, 168'h00bd6c4228e87960000001728c26273f36d7ace6af},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4148e9ba110487844c41c6a990ce6029fbacd7da, 168'h00abf5a94d89ac5ad633a85b6879affc41860f2ac5, 32'h7ffffffd, 160'h114743cb00000000000021ccc0e671308267fdb2},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{339, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6f690efb076a7dda2a0f990736ba6cd208144f1b, 168'h00abfccb16e59dd7aecddb51f4e4d2bfc2ae172f0a, 32'h7ffffffd, 160'h67063e7063e7063e7064b08f5189b9de97b88155},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=32b(4B), s=160b(20B)
  '{340, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0084b25a24491ce040eb6dc900f8ee90c6684ac8e5, 168'h0095a985e609ce016a897b913c5dff35776ceb682a, 32'h7ffffffd, 168'h00b8e38e38e38e38e38e3a4d3bd063c5600b1bb53f},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0096d267106dd68444ae300966bac62e18238042d4, 160'h5111e87654afbbad4272a264a6ba5a3320eedc2b, 32'h7ffffffd, 160'h55555555555555555555fc42fdb7e4f118d1b61e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=160b(20B)
  '{342, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c06afc4b760ec9b2dca49a4b3617e7237657191f, 168'h00f0b5ec38b9180e7ee4aa86fa19384dd28e342a9c, 32'h7ffffffd, 168'h0080000000000000000000fa647c93d769a53a912d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32b(4B), s=168b(21B)
  '{343, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0093df7994eab8a87973e7e216df0672a82114ae2c, 160'h6aa28ee71bf4154d04aed59a392761c3d1dc411b, 32'h7ffffffd, 168'h00f3574ed57ab7c5c1c0aeb155eca538ef150d0a40},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32b(4B), s=168b(21B)
  '{344, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h59ea346ba437153d58a8795b7e078689251d5423, 168'h00f113b9caa5855a8ebe9a6d0b1acf280e342a93da, 168'h0089499f94eae245d5a9b5374975ece521d855975a, 168'h00b1218927935126f18c8f57445bc5ea2a9b62ffcc},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{345, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h59ea346ba437153d58a8795b7e078689251d5423, 160'h0eec46355a7aa571416592f4e530d7f14bd56c25, 168'h0089499f94eae245d5a9b5374975ece521d855975a, 168'h00b1218927935126f18c8f57445bc5ea2a9b62ffcc},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{346, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c1329e5abc05dc8cb22c6c5e900c119fe700880b, 168'h0089643fbd2f156366b3a44316c8bb10e46e305055, 8'h01, 160'h55555555555555555555fc42fdb7e4f1437c60c7},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{347, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h1195e142718809c541296eac4d6201af46695d5d, 160'h233f099afd1ff16acb1071b4199e61e2a9c346eb, 168'h020000000000000000000000000000000000000000, 160'h33333333333333333333975b6507efc3f54aa077},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{348, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c9f7e7bc377bffc4e2a79e4836e61ed5c775dabe, 160'h073a1e62494b22fa27642f51d6f4c5d35d70db5a, 160'h55555555555555555555fc42fdb7e4f1437c60c7, 160'h33333333333333333333975b6507efc3f54aa077},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2102b319abe9060e9d4520b0b6a8ab9641b3b5d3, 160'h2b4067358970714a0f24ae1f351884a7d8588042, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h55555555555555555555fc42fdb7e4f1437c60c7},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a185a284dc8e55e796e084ca5f4ddf5bb8d70a0b, 168'h00d39ec502b4b767c9697963ec98bcd6d613c135e8, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0091c7b4456a9ec11f893316f05e8e81a7b434859a, 160'h0124d84d6dfd221aa928d768f533219eb6d5bccc, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 168'h00ccccccccccccccccccce5d6d941fbf0fd52a81df},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4549f25af5fc3a560c62f91fd555f922df271103, 160'h42890b6465457119a56148c7637a21144cac650b, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h33333333333333333333975b6507efc3f54aa078},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h7f49ac03c66731929b4ef03c7445b386d64025ea, 160'h02461eb07d492bc8afca10d37f469b14dd2d9449, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 168'h00db6db6db6db6db6db6dd1af567d8defead88f8dd},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h179d0a5fa8be0b89d8efd25948e8624e3eb1b8a0, 168'h00f614fbdda7c63019c4ad480b01a6f38b7d173138, 160'h02f997f33c5ed04c55d3edf8675d3e92e8f46686, 160'h0eb00091546e2d1fc7dcc249da653f08707af318},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00aa5cb12acdf9a8336864190c1dd6df86f98f4c4f, 168'h00b2ffdde9e2b9b558c9bfdf7aa9c7f7ec090c61d2, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h55555555555555555555fc42fdb7e4f1437c60c7},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4f052d5ded4b999f95025401553e1cd6a3f47d6b, 160'h4b4c60ab8e9ab5a0fb004224047396052236b818, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3a53aa2df4ec5bc2748e4370e608ebdd6a256666, 160'h0fdf61b9eaf36bac285002e1bfcc62e9e55171db, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 168'h00ccccccccccccccccccce5d6d941fbf0fd52a81df},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h747c6174595d49f17bb3a36c8b7166421fff8f9f, 160'h5d9784617bdd66817754e964a1c622c40cfdab3c, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h33333333333333333333975b6507efc3f54aa078},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h02489c58f2679bd170cb48776c5c6b2c6c851023, 160'h3244ffe4760912f715c443133a384ecde72e6844, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 168'h00db6db6db6db6db6db6dd1af567d8defead88f8dd},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4d0bdafb33dfb43af69e8e130dd901d129ac427a, 160'h1f74bde4f32ad5bb21ae7cae079c9fc583fe196d, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h0eb00091546e2d1fc7dcc249da653f08707af318},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{361, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h23a628553168947d59dcc912042351377ac5fb32, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{362, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 160'h23a628553168947d59dcc912042351377ac5fb32, 168'h00894b5a17a0c6db3c257d25a6ca0a19e1947c7528, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{363, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 168'h00dc59d7aace976b82a62336edfbdcaec8053a04cd, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{364, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4a96b5688ef573284664698968c38bb913cbfc82, 168'h00dc59d7aace976b82a62336edfbdcaec8053a04cd, 168'h00894b5a17a0c6db3c257d25a6ca0a19e1947c7528, 160'h24924924924924924924d9d3914ecfd51cec297a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{365, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 168'h00b0046a56f874d30ea2ba7ac1a935fd9d754ee641, 160'h7b9a54d275806819ec30b15618f5625115241f46, 160'h49c9656cd8cbee4456548d63a7fc480791909c42, 160'h6ff78980793ee086a2e66e01a490bdfc03f2d302},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{366, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 168'h00b0046a56f874d30ea2ba7ac1a935fd9d754ee641, 160'h7b9a54d275806819ec30b15618f5625115241f46, 160'h0f5720c6bd95624b603b2be5a75e487b34268d5f, 168'h00bfd6d370b516687113b12a4fc95eebb874a646fa},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{367, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b0046a56f874d30ea2ba7ac1a935fd9d754ee641, 160'h7b9a54d275806819ec30b15618f5625115241f46, 160'h2dfc21da5c39d441fc6683e54da009f413a0ff87, 160'h647382b3e39a8ac8cbe02f4666d045928a0eb061},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{368, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 168'h00b0046a56f874d30ea2ba7ac1a935fd9d754ee641, 160'h7b9a54d275806819ec30b15618f5625115241f46, 160'h4f71014057dde59269ba089c49082dab3ffa9af3, 168'h008d1abb842b2f932a04c2dd19a2f2109a57c88c32}  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
};
`endif // WYCHERPROOF_SECP160R1_SHA256_SV
