`ifndef WYCHERPROOF_SECP384R1_SHA384_SV
`define WYCHERPROOF_SECP384R1_SHA384_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp384r1_sha384;

localparam int TEST_VECTORS_SECP384R1_SHA384_NUM = 276;

ecdsa_vector_secp384r1_sha384 test_vectors_secp384r1_sha384 [] = '{
  '{1, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 384'h1840da9fc1d2f8f8900cf485d5413b8c2574ee3a8d4ca03995ca30240e09513805bf6209b58ac7aa9cff54eecd82b9f1},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{2, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 384'he7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{3, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{93, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 400'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d70000, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=400b(50B), s=392b(49B)
  '{94, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 408'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f820000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=408b(51B)
  '{98, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 400'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d70500, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=400b(50B), s=392b(49B)
  '{99, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 408'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f820500},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=408b(51B)
  '{114, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 0, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=0b(0B), s=392b(49B)
  '{115, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 0},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=0b(0B)
  '{118, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h10b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{119, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h02e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{120, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c54857, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{121, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f02},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{122, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 376'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=376b(47B), s=392b(49B)
  '{123, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 376'hb30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=376b(47B), s=392b(49B)
  '{124, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 384'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{125, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'hff12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{126, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 400'hff00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=400b(50B)
  '{129, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{130, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=8b(1B)
  '{131, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h0112b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19a25617aad7485e6312a8589714f647acf7a94cffbe8a724a, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{132, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'hff12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe1a138f7ca6eeda02a462743d328394f8b71dd11a2a25001f64, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{133, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hed4cf541094ab8901949ed51aa83fbda99e1d94bb4e401e6250d35d71ceecf7c4571b51b33ba5fcdf542cc6b0e3ab729, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{134, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ed4cf541094ab8901949ed51aa83fbda99e1d94bb4e401e5ec7083591125fd5b9d8bc2cd7c6b0748e22ee5d5daffe09c, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{135, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'hfeed4cf541094ab8901949ed51aa83fbda99e1d94bb4e401e65da9e85528b7a19ced57a768eb09b8530856b30041758db6, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{136, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h0112b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{137, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ed4cf541094ab8901949ed51aa83fbda99e1d94bb4e401e6250d35d71ceecf7c4571b51b33ba5fcdf542cc6b0e3ab729, 392'h00e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{138, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h01e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc5f8fc6adfda650a86aa74b95adbd6874b3cd8dde6cc0798f5},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{139, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 384'he7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc66a35cfdbf1f6aec7fa409df64a7538556300ab11327d460f},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{140, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'hff1840da9fc1d2f8f8900cf485d5413b8c2574ee3a8d4ca039ce66e2a219d22358ada554576cda202fb0133b8400bd907e},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{141, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'hfe1840da9fc1d2f8f8900cf485d5413b8c2574ee3a8d4ca03a07039520259af579558b46a5242978b4c327221933f8670b},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{142, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 392'h01e7bf25603e2d07076ff30b7a2abec473da8b11c572b35fc631991d5de62ddca7525aaba89325dfd04fecc47bff426f82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{143, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h12b30abef6b5476fe6b612ae557c0425661e26b44b1bfe19daf2ca28e3113083ba8e4ae4cc45a0320abd3394f1c548d7, 384'h1840da9fc1d2f8f8900cf485d5413b8c2574ee3a8d4ca039ce66e2a219d22358ada554576cda202fb0133b8400bd907e},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{144, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{148, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{149, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{150, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{151, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h00, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{154, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{158, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{159, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{160, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{161, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'h01, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{164, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{168, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{169, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{170, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{171, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 8'hff, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=392b(49B)
  '{174, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{175, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{176, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{177, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{178, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{179, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{180, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{181, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{184, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{185, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{186, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{187, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{188, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{189, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{190, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{191, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{194, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{195, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{196, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{197, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{198, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{199, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{200, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{201, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{204, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{205, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{206, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{207, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{208, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{209, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{210, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{211, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{214, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 8'h00},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{215, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{216, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 8'hff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=8b(1B)
  '{217, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{218, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{219, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{220, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{221, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{230, 1'b1, 384'h1ea4d7e33dd2cad2b412822fb60c29b7280cae718af25c51f907eb101cca981ac86a9d1a9186a1b630fb6e7079385911, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ac042e13ab83394692019170707bc21dd3d7b8d233d11b651757085bdd5767eabbb85322984f14437335de0cdf565684, 392'h00bd770d3ee4beadbabe7ca46e8c4702783435228d46e2dd360e322fe61c86926fa49c8116ec940f72ac8c30d9beb3e12f},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{231, 1'b1, 384'h00000000505a3d306890ad438d155166987fcd0d78a44fa79272ef4dcade39c852dcd5a4b23075d7651bb5c57629f198, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d3298a0193c4316b34e3833ff764a82cff4ef57b5dd79ed6237b51ff76ceab13bf92131f41030515b7e012d2ba857830, 392'h00bfc7518d2ad20ed5f58f3be79720f1866f7a23b3bd1bf913d3916819d008497a071046311d3c2fd05fc284c964a39617},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{232, 1'b1, 384'hfc000000009322da48a8586f26f148003932f6d4c0d1ce3a21798f7b651dab7642188c9061a66dc9b190e00b0290e264, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00e14f41a5fc83aa4725a9ea60ab5b0b9de27f519af4b557a601f1fee0243f8eee5180f8c531414f3473f4457430cb7a26, 384'h1047ed2bf1f98e3ce93e8fdbdc63cc79f238998fee74e1bb6cd708694950bbffe3945066064da043f04d7083d0a596ec},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{233, 1'b1, 384'h76ec0000000091b9f8b1eafd062de52093243e4eba77f18c415c92cd757f7041715e5946a839457a6b05d15758bf5c8d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00b7c8b5cf631a96ad908d6a8c8d0e0a35fcc22a5a36050230b665932764ae45bd84cb87ebba8e444abd89e4483fc9c4a8, 392'h00a11636c095aa9bc69cf24b50a0a9e5377d0ffbba4fab5433159f006ab4563d55e918493020a19691574e4d1e66e3975e},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{234, 1'b1, 384'h7d383000000000c8e8c1505bdecd51dcb34bf8a0ad3ace53a07eff629b9aeb6792a9b7fd55849e57300e24cb83cfd41d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h4a7df2df6a32d59b6bfed54f032c3d6f3acd3ac4063704099cd162ab3908e8eeba4e973ee75b5e285dd572062338fe58, 384'h35365be327e2463dc759951c5c0be5e3d094cb706912fdf7d26b15d4a5c42ffebeca5ae73a1823f5e65d571b4ccf1a82},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{235, 1'b1, 384'h3b0f107e00000000c33f3c4431329dc9f62a724c34d1f01d3b3520b01647570625a5d84e7f7770d88ad6b3f195324d65, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h009ad363a1bbc67c57c82a378e988cc083cc91f8b32739ec647c0cb348fb5c86472015131a7d9083bf4740af3351755195, 392'h00d310dc1509f8c00281efe571768d488027ea760fe32971f6cb7b57cdf90621b7d0086e26443d3761df7aa3a4eccc6c58},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{236, 1'b1, 384'h72849c623b00000000164206feda0efddeb0539b431bccd2cf1d74b25811c5abf705bb56d6b9a1be3132986a6356934c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h0095078af5c2ac230239557f5fcee2e712a7034e95437a9b34c1692a81270edcf8ddd5aba1138a42012663e5f81c9beae2, 384'h40ee510a0cceb8518ad4f618599164da0f3ba75eceeac216216ec62bcceae8dc98b5e35b2e7ed47c4b8ebacfe84a74e6},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{237, 1'b1, 384'h5310794f0cdc00000000f5976a5246e50af0aeb336f71f55f2db9a239ca36619091fbdf17a9ea99057f9fa6282c87b97, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00a538076362043de54864464c14a6c1c3a478443726c1309a36b9e9ea1592b40c3f3f90d195bd298004a71e8f285e093a, 392'h00d74f97ef38468515a8c927a450275c14dc16ddbdd92b3a5cae804be20d29c682129247d2e01d37dabe38ffb74808a8b7},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{238, 1'b1, 384'hcc968637c615b400000000ddd043d9ba734fa5ba9255ccad39c0aa38cc7cb12ce310855c71bcfa238bfb0f22969f0d30, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00bbe835113f8ea4dc469f0283af6603f3d7a3a222b3ab5a93db56007ef2dc07c97988fc7b8b833057fa3fbf97413b6c15, 384'h737c316320b61002c2acb184d82e60e46bd2129a9bbf563c80da423121c161decd363518b260aaacf3734c1ef9faa925},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{239, 1'b1, 384'ha82bcb45d5a2d583000000003c39b1cfcbe18638eb31d348344391d2a5f0aa4047c7131451d62f158e4ff8a2be60ae2f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h679c3640ad8ffe9577d9b59b18ff5598dbfe61122bbab8238d268907c989cd94dc7f601d17486af93f6d18624aa524a3, 392'h00e84dd195502bdcdd77b7f51d8c1ea789006905844a0e185474af1a583bab564ee23be0bc49500390dceb3d3948f06730},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{240, 1'b1, 384'h07a7099d24245ea53600000000058ebe28e0821ed103fdb1980c9d6ab839722ef4eeda9677fbb0f5498da96b4518756e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f6f1afe6febce799cc9b754279f2499f3825c3e789accef46d3f068e2b6781fd50669e80c3c7293a5c0c0af48e068e35, 392'h00f59cc8c2222ed63b4553f8149ebecc43b866719b294ef0832a12b3e3dbc825eeab68b5779625b10ae5541412ec295354},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{241, 1'b1, 384'h7e168cf9539beb95be11a000000000be07c6e0bdfeb58307d309cd05ad4d1144ca4be88458b9029a7a309ad3dd544958, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f46496f6d473f3c091a68aaa3749220c840061cd4f888613ccfeac0aa0411b451edbd4facbe38d2dd9d6d0d0d255ed34, 384'h00c3a74fa6666f58c4798f30c3779813e5c6d08ac31a792c2d0f9cb708733f26ad6bf3b1e46815ae536aa151680bdee2},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{242, 1'b1, 384'h5482408d92e7b7b805dbdabf00000000bd35f5ad31458f62adbe67ad0e7f7672e5c33fff10ae4bbd3c76a44dd360bcc2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00df8b8e4cb1bc4ec69cb1472fa5a81c36642ed47fc6ce560033c4f7cb0bc8459b5788e34caa7d96e6071188e449f0207a, 392'h008b8ee0177962a489938f3feffae55729d9d446fe438c7cb91ea5f632c80aa72a43b9b04e6de7ff34f76f4425107fd697},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{243, 1'b1, 384'h73058e2e9c60ed128fa60cb412000000001f383491b30e7d145935a43309d930bb03428d7ad85ce3f3b7f0e97ced1b7a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h008bb6a8ecdc8b483ad7b9c94bb39f63b5fc1378efe8c0204a74631dded7159643821419af33863b0414bd87ecf73ba3fb, 392'h008928449f2d6db2b2c65d44d98beb77eeadcbda83ff33e57eb183e1fc29ad86f0ba29ee66e750e8170ccc434cf70ae199},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{244, 1'b1, 384'hd2369784531e708cbea8be46e007000000007a1386f05819191228f18e40a35351132cb18f784a009886cfbddba23961, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00e3832877c80c4ed439d8eadcf615c0286ff54943e3ae2f66a3b9f886245fea470e6d5812cef80c23e4f568d0215a3bfc, 384'h3177a7dbf0ab8f8f5fc1d01b19d6a5e89642899f369dfe213b7cc55d8eaf21dd2885efce52b5959c1f06b7cac5773e5b},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{245, 1'b1, 384'h19a517f8670cae839c2cc49f52dadf00000000938a4514a0be4e49f25d2746de5b2af86ed089cacccae74f137dbd7f6d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6275738f0880023286a9b6f28ea0a9779e8d644c3dec48293c64f1566b34e15c7119bd9d02fa2357774cabc9e53ef7e6, 392'h00d2f0a52b1016082bd5517609ee81c0764dc38a8f32d9a5074e717ee1d832f9ea0e4c6b100b1fd5e7f4bc7468c79d3933},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{246, 1'b1, 384'h75d6dd22470f07ff7e8ee31f4c52ceec000000000c00f7cb9b77e3eb6b7fa3abfb1bd4f74df594f0a0d35de24ab25f6b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d316fe5168cf13753c8c3bbef83869a6703dc0d5afa82af49c88ff3555660f57919a6f36e84451c3e8e5783e3b83fe3b, 392'h00995f08c8fec7cd82ce27e7509393f5a3803a48fe255fcb160321c6e1890eb36e37bcda158f0fa6899e7d107e52de8c3c},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{247, 1'b1, 384'hadd32288a9999a1bcc2a60ebb1a81bf76c0000000061572f564378f31ce84dba31359b336f9597b745b8d0298df06b77, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0b13b8fd10fa7b42169137588ad3f557539a4e9206f3a1f1fe9202b0690defded2be18147f5b2da9285c0e7349735ea3, 384'h0478ad317b22a247bf9334719b4c8ee84acf134515db77e6141c75d08961e1e51eaca29836744103de0f6a4c798d3eeb},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{248, 1'b1, 384'h658f165273041c07b8b2698203febbcb693500000000046259dc5bed17be79304fa9ae62170d2eeebfa602f6a0176d31, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h15804429bcb5277d4f0af73bd54c8a177499a7b64f18afc566c3ce7096bdc6c275e38548edcfa0b78dd7f57b6f393e49, 392'h00d5951f243e65b82ba5c0c7552d33b11f1e90fde0c3fd014aac1bb27db2aaf09b667c8b247c4cdd5b0723fba83b4f999e},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{249, 1'b1, 384'h6f6c8c2d15f8c71ab1bdfd0c76eced65ce8dc6000000002d9db18077477d95303a4cbe449d3c823545d301ecd721219b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h359247c95776bb17492b7bf827f5f330fa9f9de7cc10441a1479c81776ce36cdc6a13c5f5149c4e39147a196bb02ed34, 392'h00f6ed9252a73de48516f4eabab6368fbff6875128af4e1226d54db558bd76eec369cc9b285bc196d512e531f84864d33f},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{250, 1'b1, 384'hd80da84c81a082c962cf2d39d9d29e73cec400510000000088e9fb897376e222d8bdaa59e10057b4465fbfacb8ce75e1, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00a557d1f63a2094f683429ecb35a6533bac897682775c0051e111eed6e076c48867cae005c5e0803800b050311e381cd6, 384'h2a2f871efcf03cf1c8f509e076aaa2a76f1ea78d1c64804ea5b063b0324b8e98eb5825d04370106020ee15805dbedf81},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{251, 1'b1, 384'h58d56a6e9f5c44677f46218cecf14ac83d3b7291ba000000004b5871100b047f957ffa837ca9ff1538cd20aa226af5bd, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f22bf91169b4aec84ca84041cb826f7dfc6f33d973f3c72433b8a0ca203aac93f7eed62be9bea01706402d5b5d3b0e65, 384'h7841d3bc34aa47e813a55c25203c5ec2342d838d5b4638c2705dcf4bac9c24f765b5d4c28fa3c7fda7a38ed5048c7de3},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{252, 1'b1, 384'hf4af84ea49c645fb9b6d82521d1bdcdbb4e6006b9dc6000000009fd001c4fe4115387d9960801ed27510ff2404088c3d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h009c196e39a2d61a3c2565f5932f357e242892737e9adfc86c6609f291e5e6fdbb23029ff915a032b0c5390ba9d15f203e, 392'h00d721e28e5269d7813e8a9aed53a37e652fec1560ca61f28f55ab4c262cc6214eee8d3c4c2ba9d1ba0ba19e5e3c7484a7},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{253, 1'b1, 384'h0e3bdb68603cf26a71b721be3186676a718402fcca5c3500000000eff7e3ab0511ca1ac9bf296241a91bf4fe654d6704, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h008ba1e9dec14d300b0e250ea0bcd4419c3d9559622cc7b8375bd73f7d70133242e3d5bf70bc782808734654bacd12daea, 392'h00d893d3970f72ccab35555ae91ebcfed3c5bfc5d39181071bc06ba382587a695e02ed482f1a74fe309a399eaee5f5bc52},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{254, 1'b1, 384'h5447eef2a0fc916120854ab8738c97cc2bb7edf244939d1c000000005f2224ccfabaa3ff603e62e0da05e25362d58ef0, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2f521d9d83e1bff8d25255a9bdca90e15d78a8c9ea7885b884024a40de9a315bed7f746b5da4ce96b070208e9ae0cfa5, 384'h4185c6f4225b8c255a4d31abb5c9b6c686a6ee50a8eb7103aaef90245a4722fc8996f266f262109c3b5957ba73289a20},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{255, 1'b1, 384'hb1b84a290f18a916a01327114097cd286357b9da079b2fd627000000007d6121ce46dc5a526d6f3742c22d65b486165e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d4900f54c1bc841d38eb2f13e0bafbb12b5667393b07102db90639744f54d78960b344c8fbfbf3540b38d00278e177aa, 384'h3a16eff0399700009b6949f3f506c543495bf8e0f3a34feb8edd63648747b531adc4e75398e4da8083b88b34c2fb97a8},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{256, 1'b1, 384'h304411f089bc2fc9952de809857d792f9d0f2003f004b923499a000000009bd7878d036a12c37cfef0b5fc092137eb08, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00c0169e2b8b97eeb0650e27653f2e473b97a06e1e888b07c1018c730cabfdeeec4a626c3edee0767d44e8ed07080c2ac4, 384'h13f46475f955f9701928067e3982d4ba5a58a379a66f91b74fad9ac8aee30086be6f41c9c2d8fb80e0924dedbe67e968},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{257, 1'b1, 384'h654b56eca2f5cf64f5872d1632d0fffddd00ea328adea953f047fc0000000089487f48cd08f1ae0a42fdfe10a3ad5410, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2e868871ea8b27a8a746882152051f2b146af4ac9d8473b4b6852f80a1d0c7cab57489aa43f89024388aec0605b02637, 384'h6d8c89eed8a5a6252c5cead1c55391c6743d881609e3db24d70ead80a663570020798fbf41d4c624fcb1ce36c536fe38},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{258, 1'b1, 384'h00d663434dc8a7e9afe6f5874de9af85953ae9885ee2b635f2d6d9e64200000000dd8d01527d2820994d9d0728ed1027, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00abe6a51179ee87c957805ecad5ccebca30c6e3a3e6dbe4eb4d130b71df2bf590b9d67c8f49e81bf90ce0909d3c2dab4c, 384'h7110582fab495b21bd9dda064fbd7acc09d0544dcf7699be35ad16207ffa10e8904f9241a709487ba2ba7e34430b81c3},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{259, 1'b1, 384'he37d9ed3e72fedc0879e4ea9921eb2adfc4cf344bbf4574ec5df3ab15b4a0000000087ea8cf048f97f906b501e699eab, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h50252c19e60e4120b7c28b2c2e0a588e5d107518cd61e5c7999c6d465ea134f752322d8b83f5988fcdc62bd9adb36ccd, 384'h193899352491dabfe4fc942e14ddacb200673729d61602cc0baf5732d262f36e5279865a810ce2f977f57686a0d0137a},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{260, 1'b1, 384'h515faa7acd3e17f51542deeb40e22d7ae5ab734077e3de8ba8690efb7f55650000000028e356367f6499b0761f19fed4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00eb725fdd539d7de8ea02fac8db6ec464f40c272a63e6b2718c4e0266bf1235dae330f747a6052f4319ecbe7bdade9bd0, 392'h00ae84507648ba2d1944bb67722ccd2cb94b92b59e89a1ae698c668bb57f481c42b216c23da4b1d8c0e502ef97fda05ad0},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{261, 1'b1, 384'hd4f4add5532fda6aad489da3efeff9af174e579294e8e782810d6908a25368a300000000323ea656e24f56ed7182e776, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h25aa56fcbd92f2cf53bddbaa0db537de5843290731c1dd78036fcbded4a8f7187ddfed9f5ca9d98ea7b12d24b8d29d57, 384'h028f68372d66164810bf79c30a191116d496fe32314605dc1668289425fb3a15d7532dde1052a49a35866c147abde1d9},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{262, 1'b1, 384'hfc21130bb192b7238670db30a3e1033919bb4be067cf2b2fb43a06ac794055197300000000bd0faf1c48fefa7a25b156, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h54bf7adc8548e7cae270e7b097f16b5e315158d21b0e652ce1cfe4b33126ba4a65bf227b4cddcaf22d33d82478937b20, 392'h00bfc1b8f1d02846a42f31e1bd10ba334065459f712a3bbc76005d6c6488889f88c0983f4834d0bf2249dbf0a6db760701},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{263, 1'b1, 384'h770cba8761c32c733b1065eb678fd6609273d42ec0c0da9cecc0e1a4f291961d83df00000000f920643dad519cd2544b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d3bb29ac0bd1f6058a5197f766d6ea3216c572ded62af46318c8c7f9547bb246553654279d69989d9af5ef4ccacf64da, 392'h00e10281122c2112a2a5a9d87ac58f64fb07c996a2d09292119e8f24d5499b2e8524ebd0570097f6cc7f9c26094a35c857},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{264, 1'b1, 384'h1701e1cfd87a9b14aa68513d0470d17c59efe08e7a47061ec7376249b2cd919fdfeab700000000020fdc71a9808bdd90, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00bc32e85e3112472408f9324586e525325128a38313c34b79700cb0a3f7262a90a1fcc40eef1f1a3884032a7a21810e0a, 392'h00c02f52541360358107a13dbea31f83d80397710901734b7adb78b1fc904454a28a378514ccef80ecc70c1d8e55f11311},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{265, 1'b1, 384'hd03bae59eeabef3e55e7b232af339a7e6c4b2c036f0e4702ba58378585f76852e55f120b000000004d90a75f9793e31d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f04b9e17c71d2d2133ea380d71b6b82c8a8e3332703e9d535b2c2bca9b0ad586d176a6049afa35edd9722edb5c33daa3, 392'h00bd44d4a6263380ca6f22e76c26d5f70f41f4d7cae7d4b9c1b8dc2ba5298d9d12408b04614e2f3796cc19c950c8c88a10},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{266, 1'b1, 384'hf4e5d615dfcd1d3a2e67d936d64abf4a4e8540a3af53a4e921e8b0e101c46b0f1fe19704ca000000002fdbd572673867, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00c8807351d8e261338e750cb9a52f4be4470b63f6f181cbe0e81d43b60824ba4be1bba42b1783897a0d72b0614018b02f, 384'h52e3a598c8be982127e961eed2b04f21c86df4ebcab0d955a7c66ec7f818898798ee75367a85022276b912c0a072bff7},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{267, 1'b1, 384'h4b8116f9272de6004f0010d1e05bdeddfdf4e16a2f32a8808c8b1c49e883b3f3c7934a5f05e4000000004792e40ec585, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6152841b6fb460546eeb4158a3e5ffa54f51aa6a208987be899b706055cd59d8ec7c01f4634254fe050e1d4ec525a173, 384'h73f0c5f13640d892c28f701428e8fbfb736b6478bbd972c8c684977556ed599a70d313e06b126080e13068d56e1c10be},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{268, 1'b1, 384'hcce4aaa4afd18d37eb0d3ec03e7813e3e2c9338f8e1830f54a75b1e5e8dd3456549901a6334676000000003cfb79452a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00842f8d2814f5b7163f4b21bd9727246e078ad1e7435dfe1bc5f9e0e7374232e686b9b98b73deab9e43b3b7f25416c2be, 392'h00852c106c412300bac3ba265990b428a26076ab3f00fd7657bbd9315fa1cd2a1230a9a60d06b7af87aa0a6cf3f48b344c},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{269, 1'b1, 384'h08ef3af646b01223ebae9d27e045c4a95f1b0dc5dd5a8048b17758e524e965e0be0dba299dbc3f55000000001320c4a8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00e13f6d638b9d4fba54aa436a945cfea66dec058fab6f026293265884457b5a86e8e927d699bc64431b71e3d41df20044, 392'h009832cd1b4177118ed247b4f31277da15f420179f45c71a237d77f599a45df68247bac3dcef0868ecd1665005c25b7c6c},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{270, 1'b1, 384'h54794e6b309d0a984f21a01a0a4d76c3f1c65309d1c7b41cd51de2246d76949061fe89cc162247deeb00000000acc7b9, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h09fff1c2e4ff8643cbfad588620c2bf7aaca5cf4242969142c7145b927bd82ed14f3ae8c6e2ce2da63b990b9f1be6d64, 384'h780c816f6c86343b008235ee986abf2136123ed247e4751e4d5467334f08e5e2ca1161254f68c3e6678e2d0b87d1cc7c},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{271, 1'b1, 384'h3a01a0bb7886a7fde9a7615ad9e1b96b20f8d5dd1ee53edac1f2b36ff3d69204026e793df840232474f900000000b395, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ffae6e7d2cea71b5a9c73cbc1285a8d252949772afe1aa27fb137740fc429c2a8c8648c9a5ba678a32f7ae7689b395ca, 392'h0089d54cd13a162c34189ff524813690e79768af8ebe794cc941dfe7fdf2cb8dd0b42519f034ea4d4f1c870046d13210e1},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{272, 1'b1, 384'h13d85cf840869a403889c8615682e06c23d0ce7a693fd528930fcafbf332667dc339a47d159dc05b9bc5bb00000000d7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00efa3c5fc3c8be1007475a2dbd46e3578bb30579445909c2445f850fb8aa60aa5b1749cc3400d8ffd81cb8832b50d27b4, 392'h00b36a08db3845b3d2ebd2c335480f12fb83f2a7351841ea3842ec62ad904b098efbf9faa7828b9c185746d9c8bd047d76},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{273, 1'b1, 384'h5917d7d41a220a46a2998b851d8ecc6664aa7f0178c54ef1d37be80aaa328e719ae213aea96b4a39534a142600000000, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f577095f7c74594aa1c69aca9bb26e0c7475ae5163058ecc074b03af89e56b12b6a72450589dacf0d7e6b172d0017a0e, 392'h00bee756a0b5d0a677bf95f98da512854f3ecb712f94570e1ad230eab17c527b6a8bcc9ae202b657a3611ecffa94ba0d54},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{274, 1'b1, 384'hffffffff2dd168b6e39fb11f2ba2385054725af0208ed33176168b54a1ed05ad3cee71fbe3c5a9fa8e88a7fd9bfdca81, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0ae7688c7de5882eb9c3172f5500015552f998fb53702c6cd4b03404d5a0510a8073db95db544808dbd76659fd20cf12, 392'h00bc610fe5f04d8909cc439615fb7e302d3d82992817647c50c1f467090a52b328cbbc0262f18ffb6fd9f3bd60013cea08},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{275, 1'b1, 384'h05ffffffff7cef4229da350633a4d9084d183ccd5e1823ec5471aac4f3b3d831ecadad964ea98247a4a4a08f46485412, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h5dc8a6d84afaaf900d78c6a91dc5e12e7d17891a52c1468253061d704b8940bef85b9fe807a0e02b56e8dd37c22fbb82, 392'h00914258de52932c4604dceb5ce7cc0a92e021edca9b819b84a9f25652f9af13f956a1139ee95c7aa7a079e3ad8317fbdb},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{276, 1'b1, 384'h6760ffffffff6807afd75769def299683c303d9d7e2bd99061950c64712da56e3434ccf7e8a7baace2866260564a8740, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00da55a6dbb845205c87c995b0bbc8444ffcba6eb1f4eb9d30f721d2dacc198fb1a8296075e68eb3d25ef596a952b8ea19, 392'h00829f671dccad6d7b0b8c4b39ff3f42597965d55c645fb880a66fe198d9344c9311f1598930392470379fa5ff43c75d04},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{277, 1'b1, 384'h6f9d1affffffff498199b47a27f336cca58d0961152497f7ceabcf0a9c60a2b3625c002f6301e658452c5b01dc6ff7a2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3730dfd0985de77decdd358a544b47f418d3fab42481530d5d514859894c6f23b729af72b44686058de29687b34b3b0c, 384'h65bdfaf0ac217a80b82eb09c9f59c5c8cfbf50a6eb979a8f5f63eab9bd38ee0938e4b23102112033b230a14ad2790e3f},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{278, 1'b1, 384'h7e9472cdffffffff5ea8f8066ee7b4c84a832482c10e714b7b6b8eb9da3ea3bf69e95bae5c0fd5b4de23bcaf2e891e2f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h55210df2124c170e259af1dafa73e66613aa18ced8eb40a7f66155d50d5f3124edfa55276de4797013177291e8afeff6, 392'h00c314d3a310a60647dad3318ed7f0405a64c3f94b5ac98e6be12208c8ad9835fa6b81a0ea59f476608634657b66e00ffd},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{279, 1'b1, 384'hd8754ed684ffffffff257c648476f3cbec756f28cb93cfdfa9d3279023f070b9c50be6cd0d3a055c54e24aaaeae1069f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f6c9897144b5d84964515eb0c8c3d0d9c6687c957887e93c29b2a21804b40307fb88bfd5cca11c95885d28867cb33a74, 384'h656bafca242290f7d7e9801b6cfd4bd1b07e8d7c6c1c59fd3d8e82e9846a1b2855c85420e4ee6ec2d97fec2161eeb243},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{280, 1'b1, 384'heb846f63a173cdffffffff901ee9ccb79478c01f53731793706b63782861f337b49dc4495fc1aa7a5865ae0ab6ba063e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00bfbcc5f343e2ab392ce6c1c02d91c00650c47136836a5d0622d476ac2b3274395721b1ab21882ed5cabed093b43b133f, 384'h043e9fc64c6108df73f9eced90f91185f83d89662f5a9d810c1824fbfd97b842f784305fd6b9c28c80d32d52b1538d12},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{281, 1'b1, 384'hbd7626c55e0af8a6ffffffff5ec425de708d538cef040125b332707455709362d61008fa5cd9f66122f95cf84cb6f02e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00b8f793ddd47e657a9081cbed1600fb22b38ad6a155f9c006ba98de1f383b4c0918ceea72253e0f869524b2369cd9bd8c, 392'h0096c452ff58f42e0853040a6d5c7e750b57dd4af06e2df8194e8d524e81ac000ee3315bbeabbf6a21f61b8904c55378d9},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{282, 1'b1, 384'h1323669aeac6cb92faffffffffa919616998cb4f3cbc033daa564f2f18120722257f877a2e615dfe35fcf7b8f6d8720b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h263ab1c93567e93b5ec4e380b0d3bb5ea1ce693c14a47afccc539aaf197f099d331ea9e26f1a0057148d46727acb6188, 384'h621db07ce94110e2be74fa953a00a8a554225b3f2c0f6c56b4ebd4db2f57ca2565ed3323fd708bb56ac6e28bfb40f2e7},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{283, 1'b1, 384'hffcde6e66a67646034cdffffffff1eef8cab9ce90796de58a9be57f8739867007c8421dbf90b0e4df092f6c08de15017, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h0096f4a2b3529c65e45a0b4c19c582dc8db635d4e74f0b81309696b23be920ba8ec553d4b370df4c59d74dd654bac6df58, 384'h1573ba1b280c735a3401d957ecd3b8908e4e0b7d80239ce042594d182faf2ddf811c9056aac4c87f4f85043766a26614},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{284, 1'b1, 384'h26aeeb0ba0595bd83b99d8ffffffff33c7871d47123d7314820e7acadd2a82506809c29d5c265adce54e00ecb7a7d405, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h0096a691b19a6294b311a438f8da345e480b1deaa1e940cfbf02177d5f08479976ea58aee31011d50b5542be188c9d63df, 392'h008f67dc9e1588aeb8be180013d41a036f9badfad9fe9340910cbf87243776f54bef7da2ebf3a7643866eb9a3b23fe59b9},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{285, 1'b1, 384'h2958e226692131467bf0383affffffff835f4dd2696f4bfa4cd9dbe1e614b43063d7e2a470ae6241b85f7857d9acb7d4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00cff27948c6d902c73d103d0802eb144dd89c1b0e3b9f9a5e498b0361dc122a0d555160d8c64d61539c1dbbd4bc18971f, 392'h00b60827488c9f16ba28378fd59b1a29c65073335a7f236131134674c62c8396f193c76f2395ddaaa4f24b69161eb69b4d},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{286, 1'b1, 384'h8ab4095fdf8572846b85a222f1ffffffffec5a9ebbabb6b08a5126c901892376e17b65c50725656afb9351b74f456baf, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00e90e22d9e535dfdfd86e098d5d6a0ae08f69d4a3ffaa39f6930bcf5f5ad02ee0d0472ae984edd9f0bbe5e7d63fd4f6ac, 392'h00e3f57b0a4629ecaa21f2d34a7a0834d57ba20f99c6e31b43c37811cc23b9957c8f3356f4462214d3c8e58745e50f23f6},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{287, 1'b1, 384'hdf0a780c590a26e5030b3a0fd714ffffffff98c9bb9236bdebbe6c7ddfc431a19b00245f506ee2a6563661db3afcfb9b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h18b70e272a98cc48e1e0af73146f0f972bbfbeb6b985feb2c4acd695a7a41b99c415be9c46aedaf3ddff67a65a89e387, 384'h47d6bcea088f622ad35d88bcf46d71827bcba2f57c36d6fb8a4bf2befdc0d4e3ef366d5966c4d076d3cfa43d6626717b},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{288, 1'b1, 384'h7b1f1bbb6f0579b1789e5b145a9230ffffffff38b026124a5a64772714d4ad773be8d352a5a31883132647fdbaf2efa4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00acfd981c55fd5286cfce173726d51c3d25f65b11b7673729a62167256774f7c894b74662a212c706e00cef096074162f, 392'h00f4d471c97797c24d96aec1de85a249ef468d6036cd712563aeb65cea4995f3ee85e769b874f09a08637a44a96084be7a},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{289, 1'b1, 384'h3e83f03fc730579755c9de07b01f9ee8ffffffffc810a2a0f2fd76abc89730db5a8df79e7a1eae66e53d50d1160b83ec, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f15fcbeea8b64dad5e8566a2c37913c82d6be9d9668df469bd0b591c3923a6e12644eaf697d466fa7cd513983d946a40, 384'h70063966801079351526999e5c5c2c5f627e4c8bc96784bcbe715fe7c7afcf69785d1c8c7ccd3725e364101638396597},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{290, 1'b1, 384'hfd4a68b42a044e0f93ee2d664e6afa56acffffffffa5e7af033f39d0f3ffe3bb2764fecaa791a63b129b57d171758333, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d995147939ae6d8f62bb57372227395839e25a0d4308b899d5f506cf9e0a01e8115b7e4b822f037ec95752bd9e892f5e, 392'h009bb4d07333e468f8482a790a2a2e650e2c42da8240ec5e402506b368122f046680cd71e0117897cce3df4a1555fc8876},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{291, 1'b1, 384'hcf6a074a6d661185516dfa36f481041823b9ffffffff9bf66159a9cc5709a4660da641c5f5881397bb222a6d293e0a3c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h43c6ce5184476f3f496afeae3cb96a3f9f038957686c93437b8266a233022371d266e904aa096c3566cb33824b88075e, 384'h680c13245a8bc560b638d26f0c5f261964130256939552d3fffb07b658355611612c268a89541055d3c2bf9e82cf4da3},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{292, 1'b1, 384'hb7c58195701f1afba5beb9c4c6e49a72c27ba930ffffffffbf1d4dc72e056731d4928fb5418aab897b086f49bf709087, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h447539941dc350767fc841083d25d9247a0807e1e22e0bb9d94f504f721981b413d521efbd75e4fe831ee26338cf3de3, 376'h395ab27ea782cee4be53e06c7616bbd41d6926b18d219d75d5979f13cba2f52101019b0ec0a41ffdbf29ef73ddba70},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=376b(47B)
  '{293, 1'b1, 384'h64386b3ed6d9094c46056229331338caa6add94cd3ffffffffb6b37bcce5e1489f6864d0beab480f2f5ad5ed792c8c05, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00a0ba8e8b979c20345e34fca98531900164a859923bd6986a9c39236a2f5de053a252997f35e5b84b0d48ba0f8d09aedd, 392'h00facd6df04358fcd95fa9018a6fc0828dfe319812ff65929c060b18ad4b9f06e7fc0addd1b695315d71c15e51dc51d719},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{294, 1'b1, 384'hd6bbe3d39f94bb4f82c6b2fd8d7ae4e0b8d83343f749ffffffffa398084ca2ce44c93b06fd132b5971d1b82d51aa75a4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00b8378390f71f0bb6663f1846daf6908f8c84f770ae740cc8054122494cf0ffa9437ab26040ca22808fb29a810b70126e, 384'h427636b929a500abc34d9f22977b81e734919afaf3ed2c91eeada7074e0c16bdc52f960eaec9db5a879c1e6414035101},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{295, 1'b1, 384'h57b62b08bc87cfd374c336e21ecb4cf1c5a2a948b83756ffffffff019bc82803f3d4b443d3a613ff7df4f5bf43487224, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00f36a9048fd94803d3d6d1b11430b90b94ef8d5d2ad89018c69473ce9cfe0d6105b3c2fb2e7555ccd25f65af8c872bdc6, 392'h0081254841e7ecbfd0d810afaaf5afd6d6c5d0542bb00cc183b1db01767120afbcc0006ddcba8db7baf65f302723dabc4d},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{296, 1'b1, 384'h4d75df3eadf4570f812580ec955cccd7f5b7531fc6f1c8dfffffffff15b0eb3d151f946c5f634cd622c28967db6b7bbf, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d8a4d96409c191baa9540bf35f1d5192f9352d7f0e14f92c0e8e1f19f559b42ed3c6b7bdb6becc56584fb5c09421e2e4, 392'h00d966ba13d4245e248eafb46f2a3df92c2037d5969c7db6dbcb0ff4b21850e16a18a29785267239886365cf721a212536},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{297, 1'b1, 384'hbaa4687d7f816122b9872bab05941c32509a3aaa6a1100e5cbffffffff01c5d7c2f18ce89a64f19427ca63e12924c4a6, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1d5d86fd48e65b0cf0b0b46062241f89cf65785dd818f93f1162771a38a15f20febc261812ecaaf6f4f2b86b3362d7eb, 384'h0c76e363de1432513cb9dad6493931381ecd25f142e61968b6f20d7b1270cb9e38a7ae54e4778aff4025eb00c6a67aef},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{298, 1'b1, 384'h14a722871b050d49a7d6b6d92620364e1cfc219ec267b3c5bd0bffffffffe366153701531c1889438010e2134d461a24, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0508eed148f061114be18e8a86188feabf76b873b36eadcca9c2c60e24a2002fe456231decf7a8f6f032c08dbe0ab5a9, 384'h694c0ad781b2341e30e1d0739ac99672064f48821a69852c7940cf1d621738199c980d56d2a0b71b3fc6011c6b2444ba},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{299, 1'b1, 384'heab35662fb1999230c15862e89d7e2e19731b7d777a4b5cffac9f9ffffffff1fec7ca65935120ac73955ce4167482e05, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h726ef88bb7947a043116c111cb519ddeda3e6ffbf724884a1b22c24409cdf2779d93ce610c8c07411c2b001399103d6d, 392'h0095dc1d65046caf0e8dad07b224798d6f7807278e737883e7c7bf0b446791d4ee144c26f710134861af4e6771d4082896},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{300, 1'b1, 384'hae162a45ac34fd3b3cb8b4aa99491f5384b145d4935b8b9faa913f31ffffffff45a0a7c28ea332fb5913b47c8f8c65da, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00eb0e8e3c639f5eba8eccd9020d0ec62d8ac73f3fddbdfa08fdb2155deb0a536923ebd55e20020cab9f8e39a43a88be11, 392'h00c796df399fc35883dd5dae6817d02d3d67a8eec6601585e5e36fd2c134eddb1447ec12b144dddc9aae28a84f22602641},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{301, 1'b1, 384'hc4757d55c0621c059444c654cd1fd6a1e7b7db3e44f99975c669cd794cffffffffdbb4db5f0d1ce777a8c255ad49e58a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00e8f8c69d0396ea900f9757736d2b19dbc2d2a8c01dccf490c8b9455bd63b34c095867e7cf3b84dc7c3c3d6b51bebf405, 384'h58152a7564eeb22a3e26597026d0cd7835725bd512245448cb5016eb48ea759809fd6949d0ee5d579643f72f908c16bb},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{302, 1'b1, 384'hf28ea71729613bd5bcca29e36eaa306d9683e6636026b373121d4f04d8b4fffffffffcfd13fd547359b70b888e590928, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h380b4e48b3ff012af7c08bf871d9f4da0c708b5494a986d3d80b1979e579d0dbee61db9bc3c04c396176410788e15a0f, 392'h00e6971c013c965a7e4df10f95620a5092fab096bd5b50828f4bc91c5e479bccf6e0daf287e7ef580fa9ea153fa1a507a2},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{303, 1'b1, 384'h6ddab4131e3f9e1ec8846f07a69183a80c57c6a272c521657d428a3172d98ffffffffffd6e2f7d3018ee90775475ab9b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h008061de12029e2b000d157a455ecf2301222f092df95b9551b78cf0ef3a64f12212b57ec7b16d2c0f258946f51cb1633a, 384'h0ac2ca6ad99b29ca29a0dc38b34443ee41020f81ed9087cef7681a00c4fe60653a572944ba37f1fe51d112bfffbdd701},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{304, 1'b1, 384'h209cb6971fea0b32ccc4c721287df2bf3e2d10900a7fcd250c292c04ef38e113ffffffff74ec9c21b4c60adf33e906c5, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00e74f2a791eeb7341cff6cc1c24f459e6c0109924f7984639ae387e3ceb58758a1bc3839dea1fc3a3799562225e70a733, 392'h00d90e4d0f47343268e56bbcb011bd4734390abc9aa1304b6253e78f5a78b6905aa6bf6a3892a4ae1a875c823ae5a83e87},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{305, 1'b1, 384'h5e9f272a6766953d68cc71ffe68852c5c2085c0a3d9df20e1495d35603bc10e18effffffffb37e08990a5d8b7d2396b4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6a1cd0ff7906be207b56862edcbc0d0bbfb26d43255c99f6ab77639f5e6103a07aa322b22ed43870d1ce6df68aa0a8c1, 384'h655558b129aa23184500bd4aab4f0355d3192e9b8860f60b05a1c29261f4486a6ae235a526339b86c05f5fac477b6723},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{306, 1'b1, 384'h081d6d1c08a27c5bd5d1022079c6fae88da30067a02e72fa5b908fe92e7c548a25afffffffff9049cd225e7c0f2aa678, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h0081111fdc5f0de65583c7a5668d26c04ee52e08dac227753132cff1741cb721e112aa793c0d5fa047faf14cb45dd13e1f, 392'h009a25cf1e6c152bc3e216e021561d194979f1c11fe17019ed7bac2c13c4010f209665e3b6f33b86641704d922b407818f},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{307, 1'b1, 384'h754098eae30eee355c45a45247e549b355a1018d257f7c06e51bb1f39833ad62b2c980ffffffff6e98c80a3bdf49ace2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h009b66d122a315095b2b66ccb97272c476a2d760e827fdea05732d634df3d066569c984dd941aad5f5dec4c2e1b7b94a00, 392'h0096c32403c85bc3d0ee87f96a600182796dce53d54d7467ae660a42b87bb70792f14650ac28a5fa47ce9ca4d3b2c25878},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{308, 1'b1, 384'h394e600d5b850dba7709f631c5213338964a7f8c1c5d10cea5253e2ded1ac3e4c7169282ffffffffe04a473853d08e25, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2bb062a002088d62a0b7338d0484fedfe2af7e20cebf6a4788264eb27cb4ebc3cc81c816e6a35722cf9b464783094cb8, 384'h46cc21b70f2133f85ab0443bebe9c6fc62c6e2ec1fd9c4ddf4a6d5f3f48eb7abf1ee7bdf6725879fd1b7daafb44f6e04},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{309, 1'b1, 384'h37bc45a4c75f4c2a3837c7142a260d898cb300068cabbebe331eead41bb6c1ad967e93c56fffffffff9e274922263511, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h33e87061ee9a82eb74d8bb4ae91606563c2e4db8b09183cc00d1119ab4f5033d287a1fc90a2348163fdf68d35006fd7f, 392'h0096db97c947ee2e96e6139d3bcbf5a43606bae1ad3ca28290fbad43b281ef115ec1b98bc581ef48094f8c1aa8e36c282a},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{310, 1'b1, 384'hda5ca26a4c99b6dd983dd30bc321711c28fb09e4b370dd51b9c1b50c8d3cbe30be2c10092fb9ffffffff1de6123963b2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h70f80b438424ba228a7d80f26e22ff6a896243c9d49c75573489ee0de58ec60efd103838143465bd8fe34672ba949617, 384'h115492bd9365b96f38747536318bffb819e7c146df3a5a7a46d6288c7fdf31cff570b22176aa398daba9073ab1e7b9bf},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{311, 1'b1, 384'h22daa42bf1bffb894b5ab27dd1f2ee31fb78b51386db5c38e03512ed6b70a2161caf8aed1e6f60ffffffffff5e446670, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00ff16ca0389ea6948f4305b434fe0aa589f880f5aa937767c31170ee8da6c1ad620c993d40ddf141b7fda37424d51b5cd, 392'h00ba0f86985dffc61d6e35a37de06918b11e431b72403161acfb8f05c469f1fcfa6e215c6f7eb5a0a5e0cc9e7be79ce18b},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{312, 1'b1, 384'hd0aefbc1e1ecc970df048094c6c1f11278b26272a641ca578ac60c9404b63f6c0ea5498d5e41c524ffffffffb2dd4333, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d60c24bee05f5198cd155ad095ffb956bbcfb66b82fc0d3755119915a62f2f923557b85ddc1d12e6a757f23042cb601b, 384'h2c4d968b5eac930b51d283b418fcff6df3a9d6d66e3812cd1bf5fde797fd203a7c439b1b381e4fe8b44e6f108764a7dd},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{313, 1'b1, 384'hbcd99674934bd49800c582b5271a55745b1e365b2ce18660edfd5e3ade2c014c48b0b8acf3d75a3a4bffffffffbfd063, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00bdf634d915a4fae7a155532ca2847c33a6babe7ef8db0af50f485db3dd2c8bffe722394583932f6eb5cd97f6db7561d9, 392'h00bb425cae2e5483174b5ed873af4329da4618c14458141850bee3c7bf1ffb3f2030159043277dacc708e9d32f63400083},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{314, 1'b1, 384'h91754b64495493e276038869f7d4059e4fd5d0e9d63410342fa2669e12c8bd0fcb76d458ca99840d24d8ffffffff5d43, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h061320a3bcebac33cf399d45d1e1e1b34f37288fe4753f4fddfd496eff427e1d26b1b91d749cc34c12f4ecef837c0e8f, 392'h00fd5cf468cda319fe06e773a190c38de6e150a321ac1c416ad875432cdb7a07134c446f13068e71a1a96e35da923974ad},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{315, 1'b1, 384'h896e2e5db3422ceb81fb40f9a65a2385c8d21e078994b181969ed575e6d110ab9364a8a8be347e508ca4b8ffffffff70, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h00d620f063d33efa859b623f6c9a92340e4cdd854ffbe3e5e01379177aee31715ce587b00bd0aea98fddf236d2fc8a7a74, 384'h671f4b7c187297dc236c61888b6d9397e97783077cc4101807d79ee62e4a53a78c4b6a3a31b03178668af894a3d8902e},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{316, 1'b1, 384'h3c38114a4d2c93c8d2501af3a310cb67bd399b2715dca6b5b3b5254fe6a19ce7a9cae839db4b5e5f022f4bc2ffffffff, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 392'h0091c556c5bddd529fe903b86afc0eb8fa1f49425b779a39114ae563bebc947e633ba4ee98948faa8940dfe2562c63e1c5, 384'h198b00079d8db072d25b0a49bc8bc36457926f3c101527528df6679f92c76f1b487e6695d4b92fe33b4ee7046a6a5df9},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{317, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h4bf4e52f958427ebb5915fb8c9595551b4d3a3fdab67badd9d6c3093f425ba43630df71f42f0eb7ceaa94d9f6448a85d, 392'h00d30331588249fd2fdc0b309ec7ed8481bc16f27800c13d7db700fc82e1b1c8545aa0c0d3b56e3bfe789fc18a916887c2, 192'h389cb27e0bc8d21fa7e5f24cb74f58851313e696333ad68b, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52970},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=192b(24B), s=392b(49B)
  '{318, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h4bf4e52f958427ebb5915fb8c9595551b4d3a3fdab67badd9d6c3093f425ba43630df71f42f0eb7ceaa94d9f6448a85d, 392'h00d30331588249fd2fdc0b309ec7ed8481bc16f27800c13d7db700fc82e1b1c8545aa0c0d3b56e3bfe789fc18a916887c2, 392'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000fffffffe, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52970},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=392b(49B)
  '{319, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h3623bb296b88f626d0f92656bf016f115b721277ccb4930739bfbd81f9c1e734630e0685d32e154e0b4a5c62e43851f6, 384'h768356b4a5764c128c7b1105e3d778a89d1e01da297ede1bc4312c2583e0bbddd21613583dd09ab895c63be479f94576, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52971},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{320, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00d516cb8ac8e4457b693d5192beeb6ce7d9a46bef48eecf3ea823286f101f98d130f5a26dc6fec23662eff07f14486fd5, 392'h008456932e74894b7f0e3bb0dfd362502b3765dd80a3177209fb221dc9b51aaf4470b245391405bef514176b13a267a720, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00d1aee55fdc2a716ba2fabcb57020b72e539bf05c7902f98e105bf83d4cc10c2a159a3cf7e01d749d2205f4da6bd8fcf1},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{321, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00a8380cd35026e13bf87be693cdb6e75a82d765b4019b529e8d277c4af6c9db27ebb5d3f86e88add9d5b61186f04c83a9, 392'h0092a187507c737325d2cc624acef3cd036bfa99e0c1518be65c88bb51f900f94123acabad81d15130d3ade7ff7e4364e1, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00b6b681dc484f4f020fd3f7e626d88edc6ded1b382ef3e143d60887b51394260832d4d8f2ef70458f9fa90e38c2e19e4f},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{322, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h554f2fd0b700a9f4568752b673d9c0d29dc96c10fe67e38c6d6d339bfafe05f970da8c3d2164e82031307a44bd322511, 384'h71312b61b59113ff0bd3b8a9a4934df262aa8096f840e9d8bffa5d7491ded87b38c496f9b9e4f0ba1089f8d3ffc88a9f, 8'h02, 8'h01},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=8b(1B), s=8b(1B)
  '{323, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h44ee3335fa77d2fb02e4bd7074f45e598a879c0fa822ec718c21dc13b83440edc4e3c10a1858423e03044c9eff22591c, 392'h00d027c49933e5510557d6b4b2c6f66fe5dcb9302a3b13fdc68048c3fcac88ba152b6a9833c87fdc6280afc5d11ab7c107, 8'h02, 8'h02},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=8b(1B), s=8b(1B)
  '{324, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00e2f87f72e3c66c73037fe77607d42ad2d9c4cc159893b4b9b8b0365d3a7766dbe8678b02e2b68f58e5a4f7681061a390, 392'h00e38f2142818542bef6b2bc3a2c4f43c95e5259d6bd5401531378c7ca125a1f6cc609d4fadfc5c9a99358ee77ff780c8d, 8'h02, 8'h03},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=8b(1B), s=8b(1B)
  '{325, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00e2f87f72e3c66c73037fe77607d42ad2d9c4cc159893b4b9b8b0365d3a7766dbe8678b02e2b68f58e5a4f7681061a390, 392'h00e38f2142818542bef6b2bc3a2c4f43c95e5259d6bd5401531378c7ca125a1f6cc609d4fadfc5c9a99358ee77ff780c8d, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52975, 8'h03},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=392b(49B), s=8b(1B)
  '{326, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h05e67c44fc0cbc9a8eb343b4d6f596c7d00cac5da8594caf45b7209397496214c42d856a015ce589bc9ba865a4fab5ab, 392'h0088a01c7b5d09efaf878fcb9102fb3875a8381af234d1c593076e452225a56f51674f347126d3009b44dcbb003a64d95f, 8'h02, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accd7fffa},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=8b(1B), s=392b(49B)
  '{327, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h0bb03fce3c01ebcf0873abd134a8682f5fb8dbffa22da674047e5c3e71e43de582ed6abb908c2e4faa5d96186278b6c1, 392'h00ba3b22123e68ccc56f17dd79ff15565706f71a0b6123c77af3cd88f0af024cc5259781516edcaf5fe990646e7b66999d, 16'h0100, 384'h489122448912244891224489122448912244891224489122347ce79bc437f4d071aaa92c7d6c882ae8734dc18cb0d553},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=16b(2B), s=384b(48B)
  '{328, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h58f246090d5e49863bc0bf2d501ff72f551c5f1c5e679eb49064fd02e221a2707326ec2d140bcc817afaad5065761566, 384'h497c823fd736882cbf78fb92b1a5589b67e8067497c710a4cbb39dee2c5431bc45cfb96c9f8454385c9f2b3ef2d3d31a, 56'h2d9b4d347952cd, 392'h00ce751512561b6f57c75342848a3ff98ccf9c3f0219b6b68d00449e6c971a85d2e2ce73554b59219d54d2083b46327351},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=56b(7B), s=392b(49B)
  '{329, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00fc6984dd6830d1485fb2581a45a791d8dca2c727c73d3d44c89f0082c1868af5ca74b4ca4ae22802640a9ebfe8c7ae12, 392'h00998d63a5b5ad1b72b899f0b132e4952aaa19d41fdeea48b1ed6b8358dd1db207fd66e01453ad40f67b836adc802d5fe8, 104'h1033e67e37b32b445580bf4efb, 384'h2ad52ad52ad52ad52ad52ad52ad52ad52ad52ad52ad52ad5215c51b320e460542f9cc38968ccdf4263684004eb79a452},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=104b(13B), s=384b(48B)
  '{330, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h1b8def5922303d647e8eb07e3bad92f924b79b769eef168e7541de1f4e0d28ae9733eb98cf8a1fb6dd52ca02c8c75b51, 392'h00c7aa4bf679d49d8114122074da8f6044a427371796a5654a6106162d5f686abb73ebd896ab08c7062687f12171fbe4a3, 16'h0100, 384'h77a172dfe37a2c53f0b92ab60f0a8f085f49dbfd930719d6f9e587ea68ae57cb49cd35a88cf8c6acec02f057a3807a5b},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=16b(2B), s=384b(48B)
  '{331, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h1734a039a88a16c2ff4aa97d2399121f56f52ef01ed5e50887f736f65b6e51d6e8786abb4e063da5d1ba812dff998403, 392'h00ccd698e6c296d5cd69178f8a82481a865da331627f1c4b324fbc02b36e8b5ed58a31f728e904d203a388755302195765, 104'h062522bbd3ecbe7c39e93e7c24, 384'h77a172dfe37a2c53f0b92ab60f0a8f085f49dbfd930719d6f9e587ea68ae57cb49cd35a88cf8c6acec02f057a3807a5b},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=104b(13B), s=384b(48B)
  '{332, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h52ca47dda99172cb8321495acf988548295988ec973c1b4ea9462c53e5768a704a936410ee847b5dbf1e9d0c131da6c7, 392'h0087a47027e6655792eb002d4228ee72f7c814c9a0cecbff267948f81c9903ac10eb35f6cb86369224ed609811cdf390f4, 392'h00ffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc528f3, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{333, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00bd3d91f003e18adbea73079d4eba23b91fc17fcec14c9eb15a193fbc9ca39c8c747cd7a2c9623e05dd587ccbb8ab4c44, 384'h3adb0a0706aa5ea7a68042082fccefc979612a7a1a3d694b00793b03f89bff866a8b97c8e77990c29360ce795036c764, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 8'h01},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=384b(48B), s=8b(1B)
  '{334, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00bd3d91f003e18adbea73079d4eba23b91fc17fcec14c9eb15a193fbc9ca39c8c747cd7a2c9623e05dd587ccbb8ab4c44, 384'h3adb0a0706aa5ea7a68042082fccefc979612a7a1a3d694b00793b03f89bff866a8b97c8e77990c29360ce795036c764, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 8'h00},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=384b(48B), s=8b(1B)
  '{335, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00f896353cc3a8afdd543ec3aef062ca97bc32ed1724ea38b940b8c0ea0e23b34187afbe70daf8dbaa5b511557e5d2bdda, 392'h00c4bd265da67ceeafca636f6f4c0472f22a9d02e2289184f73bbb700ae8fc921eff4920f290bfcb49fbb232cc13a21028, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{336, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h370d9e2e31c712c8028092f802319d7fdf5b3319a8518d08bed3891508c7060cfe2236e18fa14fe077093ceae633e543, 384'h0fd79aacf9d16ecc19b12d60fba4998dfc682702ec7c8bdd4a590035773b8c9c570ac7dcd414e03252f7a0e6f53b5863, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{337, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00941e6cfa356e572dcccaeb594b06955d99dc4bf07958fc98ffa17de11c7521bf2c7aa8ff260952fcb7aac078ede67b47, 392'h0090a78a0296b041a10f003df1998da4cc4a1614ebcbf5d239431f33d90d3023edc1802e8db6dabcbae67cc314da2aabab, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294ba},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{338, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h3ecfd58a3ce583866e0471d16eb3c10a411ec3b8671f3a04769b1ed8464a71cf1c76d8d9b7e3670bbe712d6f554a9383, 392'h00d980d8bedf57470d6b45cc1ad0c6426dc70a0e4be901106a36663bfcab04fcb86008777b92445120d5e3641d97396362, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 392'h00f9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{339, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h4150ccd0fa45aa2ef6b5042ddbb1b87c5ffd1115a8fe5995641948acda82a7b190762d84352cd74d1ca01e79f68f9cb4, 392'h00eb11be9d494c181c156e23e77e532bdf0a20c3cc74ba8c29b1f3eb2bd99129ee0d70ff0d593f0d7a6d6887e7c55930d2, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h064ed80f27e1432e84845f15ece399f2cbf4fa31aa837de9b953d44413b9f5c7c7f67989d703f07abef11b6ad0373ea5},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{340, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00e78fe2c11beac7090ee0af7fed469a8ccebd3cccc4ee9fccc8ef3fc0455b69aaa082dc13e1d84f34026cb6f0af9e992f, 392'h00f34ebba71bf3a4050bf28e4084b5c5f5d4098ec46f10a31b02fb4bf20cc9362f6f02a66e802f817507535fac3ec0b099, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{341, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00ee24ab8a34d05af684939357f32759cc5a14f3c717529a20aea8e0c5965d8a41e68925f688471994b72021ba51b28c09, 384'h0a55693c92ad0cbae9edcf515e2b4c060b888d82c81e4a3b6a173b62ed04a46fa95db1a2f3949980fba2e371263c4fa9, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 392'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa84ecde56a2cf73ea3abc092185cb1a51f34810f1ddd8c64d},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{342, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h3d2e916055c92e1b36133f5937b37c1b0102834eb77008a3ba9c3da446e9065971d68ba913091851e10cff5b4cd875c1, 384'h39aa7aadfc2caf7107b17ae1aea8b299d61bf15aca0cb3fd6f1ffde8192bfe58f0822bbbc1f55bddf6b4fe9c8f2b0eac, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h533b0d50480a3ef07e7e8af8b1097759bc03ac9a1c7ed6075a052869f57f12b285613162d08ee7aab9fe54aaa984a39a},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{343, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00ae596697427aa250156c05ac4338e48980a7f093ea1f1fe67098b43f6539c1b20ae74338f9bf270d33663c50abe8fd00, 384'h1ca6a52732db74ab15d2f249a3d839080f898367dfd64992cdce2708deaad523a2a236b43400424241c91a35b530fa50, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00d49a253986bbaa8ce9c3d3808313d39c3b950a478372edc009bc0566b73be7b05dad0737e16960257cc16db6ec6c620f},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{344, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h0088738f9981dd4d1fabb60ad83c2dd6dfc9da302209ae3e53498a883b6e39a38bead9b02709f352d3e6b6578154eab252, 392'h009388a05c6b9f3a4028abb9950a51f5264ecd7580a423fdec9472faeeb57f92e31c46bef2a781fe5edad026009f198262, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h285090b0d6a6820bbba394efbee5c24a2281e825d2f6c55fb7a85b8251db00f75ab07cc993ceaf664f3c116baf34b021},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{345, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00f421541311c94fdd79fc298f8ab1a3adfd08029fdad439a94d4cea11f7e799bc439609f2fb7be3f349d55e484d0a0d36, 392'h00b35330bbdbec1e75f2984483d96bf210d722c1830292ffc35a2f6a21a4b50519f565f024bbccc97228a2f8ad8fadc0d5, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00b39af4a81ee4ae79064ed80f27e1432e84845f15ece399f2a43d2505a0a8c72c5731f4fd967420b1000e3f75502ed7b7},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{346, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h399be4cfc439f94f2421cbd34c2cd90bae53eb60ddfafca52f7275d165d14fa659b636713b5d4b39e62fd48bae141d0e, 384'h1b23e3b4f0c202ed7b59db78a35c12ac698c603eab144fd09ac2ed8f4495f607e4d2c87a23ce2ec33e410ca47ecc2555, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00af4a81ee4ae79064ed80f27e1432e84845f15ece399f2cbf28df829ccd30f5ef62ec23957b837d73fe4e156edccd4465},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{347, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h1578bbff72137c4bca33d7385a892be94cb059f9091ddfe890345f712a9fba5fc77084cec11084ed048491604a07f66c, 384'h76bbaa872f0710d82a08d9dddd833c7be7c7e8e265f49145157eb4e8e8280076a37ee5873271db510034da19da24415b, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h5e9503dc95cf20c9db01e4fc2865d0908be2bd9c733e597e8a5bb7b7a62abdff6dbe3978ae56536d0fb01172ecd55f57},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{348, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h33ba451c85e729058f83041077a4695eb47df93e718b09a4618c753ac803cd75c1a91290c2ff5a635389d07149571dab, 384'h1fc7d8a71776851ff244ff632fe6f92e1652e5284893c4244fe775d8efc589d823dd03f3919027f004537bd8ee09f3a3, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h1ee4ae79064ed80f27e1432e84845f15ece399f2cbf4fa31a3ae8edab84dc3330a39f70938e3912bd59753de5aed3088},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{349, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h040771e3390216fed2c6208bdf5bfea83ab1915b166e626569f12efd410a39b7e7c76f70f0012843a26debf4ccc33dda, 392'h00e5bc5f7e62d054eac31cd022afdb71b7c638f24c30cbad0ef35ed2fc9917f356e9c3f04391b21d1035274b81537fcbf3, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00bb51cd3ba8eb201f53ddb4e34e08c0ff7dff9378106784d798d5a3440bd6dc34be3a0eaef8776619a0c97fefb15720b3},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{350, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h0098d3f16e1c510a933e648e78d01588319f002e9475df8942a2a89db0666bb7c88b32bb248140e44ac4ab28111b2b7923, 392'h0099a926f4a66fbe28ff65c09f8306893aec094b89d0fe529e3577c5ecf30a7944caaf530f4575eb113fcf4c200d2dd4bd, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00e707e267ea635384a6da09823149f5cb7acbb29e910d2630c5fb5afbc42aa8436349b214a3b8fb9481ec999e005091f8},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{351, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00d1fd602feef80be9e55a19d1a9799c72a899110c6ac21fb3c21357069809d591a8775b64d1867a8cfff124f6a5e3a4f5, 392'h00f9548064f01b9af8868705493a37a037193b48f53b7c7973023f53e6ceff6830ca2f7a14ef51536d453af43b3058d8a9, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00acc4f2afb7f5c10f818175074ef688a643fc5365e38129f86d5e2517feb81b2cd2b8dc4f7821bfd032edc4c0234085d9},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{352, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h0082f37604f66664c2883dba6d98397c281045cbf59f1d16dddb1381126a246553a8b4d2aaea48ad9185a1645f65567d31, 392'h008a4d7b19f1d2e4434c9a8ecad396304abc82221bbab0679935071c72fd975e7b021c04b1d16ea36fc2d051ef5a8e117c, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h0083276c0793f0a19742422f8af671ccf965fa7d18d541bef4c05b90e303f891d39008439e0fda4bfad5ee9a6ace7e340c},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{353, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00f052dfc27bf8a6d36f3739f239b981f5b53fe08d999ec683b01e43e7596156206ba08b8b9f59229e2fbdce05f1e40f99, 392'h0090f0fdfb7029f9b3e8c6144dad0339208b7cdcb3820a554259db9d27afdd18f4a750296c59bad6b62df076f90d53be0d, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00942848586b534105ddd1ca77df72e1251140f412e97b62afbf85d4822309176b5965453dee3fab709e14156b3dfcecca},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{354, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00f877bd6e2a9273e322a3298ea3add13d1104b32172283669ca6688f0cb591524a7f15dd41496681eda98939aae729fed, 392'h00e85ca37c81ef19e3dc9ab16908a3720d86875a51a6a6d932e37492a6ec7a344eabc482377f14891fbd1da7faeffa1178, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffed2119d5fc12649fc808af3b6d9037d3a44eb32399970dd0},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{355, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h14249bbcfeeceab06c75654d361c0df8d56b320ea3bc1d4627ec0a2f4b8fa3577445694664f569a91f480741381e494a, 384'h28479f2186d715a56788f67073056aa0cb0b6a7f7893e77b9a6976ef6663d80226896d7f43bb502e1b4d49558a27dd8b, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h79b95c013b0472de04d8faeec3b779c39fe729ea84fb554cd091c7178c2f054eabbc62c3e1cfbac2c2e69d7aa45d9072},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{356, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h50a438c98ee94025ce13e27d36b8280d4843585836eb47011a070cd77729245684a0db31fde980620349c796832b2c6c, 392'h00bdb72dba9f3f9cc878559f50b6bd1290f10a6bccbc1eeef7708b1b72059022987979e35221c51259f337c7288a2f86bc, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00bfd40d0caa4d9d42381f3d72a25683f52b03a1ed96fb72d03f08dcb9a8bc8f23c1a459deab03bcd39396c0d1e9053c81},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{357, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h4d3fc5dcfaf741113cda3ce2f8dff4c912143e4d36314c361d7ed5656b68448bcca114ba9e8124281234660b7726ddcd, 384'h680ddfef7ea07bfbcede10803d38d7211631ca11466078819eb66e11921ab7ffa3c4560c732e77595fd408e917dd9afc, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h4c7d219db9af94ce7fffffffffffffffffffffffffffffffef15cf1058c8d8ba1e634c4122db95ec1facd4bb13ebf09a},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{358, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h63d65cdfeb1f1a42000f43bd1ddd130537a7b6f635e8d2bd81a97da168221183da433ca78429fd2b33c5f94895a9c13a, 392'h00a9d1d5ea328725653a5a9d00f85a5516236f3b1428a8629287d3b0487a2e82dd57f93bb2aa3d9783dc74131e13756034, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00d219db9af94ce7ffffffffffffffffffffffffffffffffffd189bdb6d9ef7be8504ca374756ea5b8f15e44067d209b9b},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{359, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00d22c9c348b9745711f57debac3a07df90a527c06bd02a8454f41437d54224e071698f03fdc64b1d652414edc3f2239c4, 392'h009ae9812a4b92f099d6659a659691768d57e530ed3c91d5455781605850997a58221f22a2451c3932470606c23f3ab1b8, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00a433b735f299cfffffffffffffffffffffffffffffffffffdbb02debbfa7c9f1487f3936a22ca3f6f5d06ea22d7c0dc3},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{360, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h31f05c0c29e9da49aa2fbbedee770c68d10f85e7f77e72ac3cfa9c8623a2bb42eeb2f24ac8f2aef7ab0c4b4782314003, 384'h5bb32fc1ec04bbff5eab96e070c938ba1b53fe63970f649ae02e2a4ada420a249b6f7c525e2c4b9b0d5562ae26f2278c, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00b9af94ce7fffffffffffffffffffffffffffffffffffffffd6efeefc876c9f23217b443c80637ef939e911219f96c179},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{361, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00bc26eec95e26c980bc0334264cbcfc26b897c3571c96ce9ab2a67b49bb0f26a6272fdc27806d7a4c572ae0f78149f1f3, 392'h00c8af5f41b99d2066018165513fb3b55e4255dcd0659647ed55e1e2602cae4efbd6eae1dfe2ff63e2c748d4acc7430139, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00a276276276276276276276276276276276276276276276273d7228d4f84b769be0fd57b97e4c1ebcae9a5f635e80e9df},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{362, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h6fa0964dd054250af176891c0c822b013b70f059c347172cafc6b36cd16cf3b0f9d19f2598bd0d580ac16c46acb167d4, 384'h375bef701c002dcc040fd54824b14cc2df0154eb20e74464e1fe7b833426dd7d636bf2d79603fdde5ddaab23ab0cf426, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h73333333333333333333333333333333333333333333333316e4d9f42d4eca22df403a0c578b86f0a9a93fe89995c7ed},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{363, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00baa4e712ee0786a5ab0e5a5dafdcdcf87b38830ab2ec86faedda9fdf65332f6a9688269412f050356530d4664a7fb8cd, 392'h00ecc46a901b016e6bb8a336ad9aa6f19abf9ada69705d1c905beafb95a44f52af43de4bf80c050cf996b7796dfcee8e1b, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffda4233abf824c93f90115e76db206fa7489d6647332e1ba3},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{364, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h0081e78a52ae0695583f7a601ab9b6fbfaf434f2befa1f8c833d59deb627a927c2f42d48eb617fe042f584e105c23c2317, 392'h00cf22d565f5f3b425ef7937df629b6864dac71264b288c1a987210f523071319ce3f64411910ac23765c4266e615112bc, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h3fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294bb},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{365, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h41fa8765b19d3108031e28c9a781a385c9c10b2bfd42e6437e5c4bd711cf2a031750847d17a82f9376a30ae182a6d6e7, 384'h1c20af96324147d4155a4d0c867ca8e36eba204fbed2087e0fcbdc8baabe07bb3123f9f7259e771cd9f1ad17d1a23787, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 392'h00dfea06865526cea11c0f9eb9512b41fa9581d0f6cb7db9680336151dce79de818cdf33c879da322740416d1e5ae532fa},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{366, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00e585a067d6dff37ae7f17f81583119b61291597345f107acffe237a08f4886d4fdf94fe63182e6143c99be25a7b7d86b, 384'h572c1e06dd2c7b94b873f0578fcb2b99d60e246e51245d0804edd44b32f0f000c8f8f88f1d4a65fea51dbbb4ab1e2823, 392'h00b37699e0d518a4d370dbdaaaea3788850fa03f8186d1f78fdfbae6540aa670b31c8ada0fff3e737bd69520560fe0ce60, 384'h64adb4d51a93f96bed4665de2d4e1169cc95819ec6e9333edfd5c07ca134ceef7c95957b719ae349fc439eaa49fbbe34},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{367, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00e585a067d6dff37ae7f17f81583119b61291597345f107acffe237a08f4886d4fdf94fe63182e6143c99be25a7b7d86b, 392'h00a8d3e1f922d3846b478c0fa87034d46629f1db91aedba2f7fb122bb4cd0f0ffe3707076fe2b59a015ae2444c54e1d7dc, 392'h00b37699e0d518a4d370dbdaaaea3788850fa03f8186d1f78fdfbae6540aa670b31c8ada0fff3e737bd69520560fe0ce60, 384'h64adb4d51a93f96bed4665de2d4e1169cc95819ec6e9333edfd5c07ca134ceef7c95957b719ae349fc439eaa49fbbe34},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{368, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00b4d78cccbced8065c0ebdc330b4670ec99309273e442b9be341196c1043e4441fc57b914085595bfc755c64fc409f0ba, 384'h01fee31cbbbaed5c1323f09c87df9b0712c12e99733fa23ef91b4e6ca666b09dd7540ebf1068a15155bc069e3d595c8c, 8'h01, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=8b(1B), s=384b(48B)
  '{369, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h6e3c68be53aade81ef89e096d841e2845a23331e7ec8a6a839d58d07fa016c0973ed75de4f99177bfdc74db566e9d15a, 384'h4972ea08e577ce1f61c13a6ca1bad1deef2982ee01a2826f002b769f2c46098d3baff068a405d09ca3840d2fafe4e46e, 392'h01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h33333333333333333333333333333333333333333333333327e0a919fda4a2c644d202bd41bcee4bc8fc05155c276eb0},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{370, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00b101cdb3eba20e112adbb4bbd2cb479a69e590a44ea902631832abfab8af2c3041b3df7f1665b2c6eb533f546217100a, 384'h1a61aa9951578ad4f00ae17339a8a6f1359bbd0ac355678ed4df21338f08763c1d3702ec132b634c7bcc0118efb1d0dd, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h33333333333333333333333333333333333333333333333327e0a919fda4a2c644d202bd41bcee4bc8fc05155c276eb0},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{371, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h6761044a040a4979db269b4a377e42f11b4be0ce24611f677674dcf770f5887ca4db565303283809e6d65f7fc6bc2736, 384'h05c7daa403fca53549f75ff3372909642d02b7fdcac1e68242814d6e925ab01a80836cfbb35581960079e2fb44c0d186, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{372, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h6922c591502f01046fee5617bf16496f58398822e69afa8335308f36c09a8ed437209fefcffbbdf0a4876b35a3c7ab26, 384'h55854db825b94b3f27e5f892d3bbb6c7240ec922894dd3598e91fcc6134a2b8fd154e1790466906206f0f623416e63a1, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{373, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00892dac0e700fc29d1802d9a449a6f56b2172cb1b7d881013cd3b31c0edb052f2d340c8995a4477bcb9225fec15667233, 392'h00cc6c34ae17445444516fd8fd22ee83f79eb0771ebff6677ac5d4e089f87a1c72df957acb24492adcd7c3816b8e0c75b1, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h6666666666666666666666666666666666666666666666664fc15233fb49458c89a4057a8379dc9791f80a2ab84edd61},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{374, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h01634117e6478ce0568b0a2469237bbac6ff096acb7e514072bf77123cb51ba0cc3e8d69284d534d8e6d1e876cecf222, 384'h31e5ef04dc96762ce7d5ef3348ad1e241ac797ae3b630ea249afc5139af49b8ef68b32f812d6b514210363d498efc28c, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 392'h0099999999999999999999999999999999999999999999999977a1fb4df8ede852ce760837c536cae35af40f4014764c12},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{375, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h675bdc79d8243887fe1b305d12ac10d2e9c0bde070a6e3394cd5f6adfbceda75498b0e7a794c7212f42be93f61674456, 384'h3e96d1bf6f95cdbefa774911ba06463d8a90a0c9d73c9699b061d779dc52496e8ee9b9ae9c5d4d90e89cd1157d811895, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 392'h00db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6aae76701acc1950894a89e068772d8b281eef136f8a8fef5},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=384b(48B), s=392b(49B)
  '{376, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h0fd1aab89f47b565b8160dfcc433b6408adeb1473c036b26b7ddec714fb4d0e7dd756c88469e86e218813ead8e8e7676, 392'h00f1cc955c4139e0071c0079ec1d77164e0569bdf453837e8b33c98535a0e7c9c61ef24762067bb46b6116ea7909a69b23, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h0eb10e5ab95f2f26a40700b1300fb8c3e754d5c453d9384ecce1daa38135a48a0a96c24efc2a76d00bde1d7aeedf7f6a},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{377, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h34d74ec088bab6c6323968d1f468993812f690d6edca5b97604d718e12b8cdfdd96d42e57d33afe312f0ee3c3d0a13f7, 392'h0086f4922bb2c13bdf7752a3ecb69393e997bd65461c46867ebeef6296b23f2c56df63acfde648f3f5002dbc239ffd1582, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{378, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h4376c9893e9277296c766a83abbe36b34da7a631f8cbfd32a1888de0dd1455a21a153ea2d61cfa5071fc6be12a658f6b, 384'h290ba1a8ee8c78b5dd58f9ffcacb22955682eea02429c3fa8cdcb649fa4d007c8693e3f8f3c0a5f3c4de7a51beaa9809, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{379, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h10878fc4807f6732a23c883e838e38c787f7088f94c1824b84673e8b9eab16de1544ae4bf2c6fe3fe4fb343b7487e2b4, 384'h3036ff439533d22f951dae966584bafb23b217dcad2f8f4e0e6999c0c4d0f076634be805f676fd2a59c27f9fe7c5d95b, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h6666666666666666666666666666666666666666666666664fc15233fb49458c89a4057a8379dc9791f80a2ab84edd61},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{380, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h036b253e3b4ac88bb8585a2b32b978766a931e5ad0d0e653a2e34b44d6ddcc0d386e20c4def2d8bb3f8da128c1eac69f, 392'h009c8e3b5ff5dde2205af359b3974d52758d7abae812b8b275e1452c4e59cb62e9b6771d347dbd1dea761c70291cc5e0a6, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 392'h0099999999999999999999999999999999999999999999999977a1fb4df8ede852ce760837c536cae35af40f4014764c12},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=392b(49B)
  '{381, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2783c1be922fce155864ecb41d0a316e193a55843e80192f1fe556772f3debd04b9fc93c27bc6f353938886a40441994, 384'h1a352cec336946424fa3c208ea7105f5549edde8688abd305344bf4f66dda7eabcda6f8557c9af88109804d702e9670b, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 392'h00db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6aae76701acc1950894a89e068772d8b281eef136f8a8fef5},  // lens: hash=384b(48B), x=384b(48B), y=384b(48B), r=392b(49B), s=392b(49B)
  '{382, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00fa92538cdc740368caf16480ff1304cebbbe59a46a7a84603726b9592d105be069df1c61b5974f27e7552f797de97cdb, 384'h620e03a46da862e4b089bafbb80df8f055c8f47991b3a3ddb2b089aedb2f15841a6a5b5e14c1dc36b3c155c4f74d3409, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h0eb10e5ab95f2f26a40700b1300fb8c3e754d5c453d9384ecce1daa38135a48a0a96c24efc2a76d00bde1d7aeedf7f6a},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{383, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h3617de4a96262c6f5d9e98bf9292dc29f8f41dbd289a147ce9da3113b5f0b8c00a60b1ce1d7e819d7a431d7c90ea0e5f, 392'h00f9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=392b(49B), s=384b(48B)
  '{384, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h3617de4a96262c6f5d9e98bf9292dc29f8f41dbd289a147ce9da3113b5f0b8c00a60b1ce1d7e819d7a431d7c90ea0e5f, 384'h064ed80f27e1432e84845f15ece399f2cbf4fa31aa837de9b953d44413b9f5c7c7f67989d703f07abef11b6ad0373ea5, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},  // lens: hash=384b(48B), x=392b(49B), y=384b(48B), r=384b(48B), s=384b(48B)
  '{385, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 392'h00c9e821b569d9d390a26167406d6d23d6070be242d765eb831625ceec4a0f473ef59f4e30e2817e6285bce2846f15f1a0, 392'h00f9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{386, 1'b0, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 392'h00aa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 392'h00c9e821b569d9d390a26167406d6d23d6070be242d765eb831625ceec4a0f473ef59f4e30e2817e6285bce2846f15f1a0, 384'h064ed80f27e1432e84845f15ece399f2cbf4fa31aa837de9b953d44413b9f5c7c7f67989d703f07abef11b6ad0373ea5, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{387, 1'b1, 384'h38b060a751ac96384cd9327eb1b1e36a21fdb71114be07434c0cc7bf63f6e1da274edebfe76f65fbd51ad2f14898b95b, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 392'h009a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h32401249714e9091f05a5e109d5c1216fdc05e98614261aa0dbd9e9cd4415dee29238afbd3b103c1e40ee5c9144aee0f, 384'h4326756fb2c4fd726360dd6479b5849478c7a9d054a833a58c1631c33b63c3441336ddf2c7fe0ed129aae6d4ddfeb753},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{388, 1'b1, 384'h5340980991c93d7111312700b83e9e61eed0977c5bca41d5dc9e26a7af4dbef3908df6661e32e039842176176609ba8f, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 392'h009a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 392'h00d7143a836608b25599a7f28dec6635494c2992ad1e2bbeecb7ef601a9c01746e710ce0d9c48accb38a79ede5b9638f34, 392'h0080f9e165e8c61035bf8aa7b5533960e46dd0e211c904a064edb6de41f797c0eae4e327612ee3f816f4157272bb4fabc9},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=392b(49B)
  '{389, 1'b1, 384'hf9b127f0d81ebcd17b7ba0ea131c660d340b05ce557c82160e0f793de07d38179023942871acb7002dfafdfffc8deace, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 392'h009a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h234503fcca578121986d96be07fbc8da5d894ed8588c6dbcdbe974b4b813b21c52d20a8928f2e2fdac14705b0705498c, 392'h00cd7b9b766b97b53d1a80fc0b760af16a11bf4a59c7c367c6c7275dfb6e18a88091eed3734bf5cf41b3dc6fecd6d3baaf},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{390, 1'b1, 384'ha5a2cb4f3870291de150e09ee864f3b2b3b342937ac719a149439185ad6a47bb4f23ae83ff20f0c8f0c79a1764244a63, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 392'h009a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h5cad9ae1565f2588f86d821c2cc1b4d0fdf874331326568f5b0e130e4e0c0ec497f8f5f564212bd2a26ecb782cf0a18d, 392'h00bf2e9d0980fbb00696673e7fbb03e1f854b9d7596b759a17bf6e6e67a95ea6c1664f82dc449ae5ea779abd99c78e6840},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{391, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00ffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 392'h00acbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'h07648b6660d01ba2520a09d298adf3b1a02c32744bd2877208f5a4162f6c984373139d800a4cdc1ffea15bce4871a0ed, 392'h0099fd367012cb9e02cde2749455e0d495c52818f3c14f6e6aad105b0925e2a7290ac4a06d9fadf4b15b578556fe332a5f},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{392, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00ffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 392'h00acbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 392'h00a049dcd96c72e4f36144a51bba30417b451a305dd01c9e30a5e04df94342617dc383f17727708e3277cd7246ca440741, 384'h3970e264d85b228bf9e9b9c4947c5dd041ea8b5bde30b93aa59fedf2c428d3e2540a54e0530688acccb83ac7b29b79a2},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{393, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00ffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 392'h00acbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'h441800ea9377c27865be000ad008eb3d7502bdd105824b26d15cf3d06452969a9d0607a915a8fe989215fc4d61af6e05, 392'h00dce29faa5137f75ad77e03918c8ee6747cc7a39b0a69f8b915654cac4cf4bfd9c87cc46ae1631b5c6baebd4fc08ff8fd},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{394, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00d1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 392'h00c6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h3244768016457c463b74f2097f216d9670b191f76281c74bc6a1a1971d19f209bf4696468f5eb75d6326a0a43c0a6529, 384'h501e0ad985ed9f95697bd17fdbe3f9ca92e0f76426d3664e6896648d9c750bf588d0ce7d011c1a1e8d6c2e082422dc93},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{395, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00d1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 392'h00c6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h5e1af40f2480e3d97c4ae4bfd34a9f45269241356f3a46becd86a4a7c9716d73ca5aebdb3db1a7765650666683bc856b, 384'h7e7c4b473a2baaa4953785be8aa2a10006f6d36b400ab981864d69cecec046718d0404b9647454b159aa5a92d76d7955},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{396, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00d1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 392'h00c6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h6688e36a26f15bdc1c3f91367f8a7667f7bb3e30a335d6f0900e9534eb88b260cb29344c723fedfbe7ac9c5a33f4bf0d, 392'h00aa35fddf0fdc9017860b378f801cd806f3e2d754cd2fd94eb7bb36a46ce828cef87e9ebbf447068e630b87fee385ad8f},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{397, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 392'h00e6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 392'h00d4a8f3b0b4d3a5769e3a0bbc644b35f1d509355ed1fe401e170f667b661f693b32598e8c143a817a958982845042bb48, 384'h04cc07578bbd1981dbf6e8a97a354c98d41b8b6f6e8a2c2b1763c7c2a29d79e24f8476075c9aed9aec6c64dff50461ae},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{398, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 392'h00e6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 392'h00c286d1928e9c79fdd3bebdf22a1dbd37c8105e8ecf41e9e3777fe341b6b8d5a89b9d986827d6d1dbb381cd8239484a22, 384'h201119ae305b9360aa9b5e5d1567e0674c09e4f025556ebf81b987466b0f421b8d31f72bbe95f3ce2aa9874a84edfd40},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{399, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 392'h00e6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 392'h00d9c678550167f10c511e62acb4bd0a3f7f336bc090c94e6c6b02622439c348a2159c5f41f9b5aa4b470590d40dcd7cc2, 384'h1fd5eaee295abb4081cb626745f4ad279ceb44604062830b58e6c0465c562d41f02ba588fc0db1ebbe339cdc008d7a1b},  // lens: hash=384b(48B), x=384b(48B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{400, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 352'h2b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 392'h00d1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'h20fee7c71b6cb0d1da3641ec6622c055a3b16a1f596c64b34da1b2d0b868b66a8f0a0d0db983b3dc7e53bb7295da8197, 392'h008141a931d3579aec1cac9887d2fff9c6f12d47a27e4aab8cf262a9d14a715bca0b2057cbc3f18b6fd3d1df76f7410f16},  // lens: hash=384b(48B), x=352b(44B), y=392b(49B), r=384b(48B), s=392b(49B)
  '{401, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 352'h2b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 392'h00d1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 392'h00913eecc559b3cf7108a65d6cc3076bfdf36c6f94dcc6693d06690470f34a2e81564241e1de5f5f51421de30af467f10f, 384'h649bd3717244e8ef3c6b0eda983f84dca5ea86d1bec15386b9c473ec43a8cd0ba558eee819f791d9ff9272b9afd59551},  // lens: hash=384b(48B), x=352b(44B), y=392b(49B), r=392b(49B), s=384b(48B)
  '{402, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 352'h2b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 392'h00d1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'h23855c46403a97b76cbb316ec3fe7e2c422b818387604bda8c3d91121b4f20179d9107c5f92dedc8b620d7db87fccccd, 384'h50f57343ab148e50662320c4161e44543c35bc992011ea5b1680b94382cf224ea0ec5da511e102f566cb67201f30a2ee},  // lens: hash=384b(48B), x=352b(44B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{403, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00fb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 352'h208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 392'h00d200958d491fcebde667cd736c9dba0961c70db2ecaf573c31dd7fa41ecca32b40b5896f9a0ddf272110e3d21e84593a, 392'h00c2ecf73943b9adce596bac14fce62495ae93825c5ff6f61c247d1d8afcba52082fc96f63a26e55bccfc3779f88cfd799},  // lens: hash=384b(48B), x=392b(49B), y=352b(44B), r=392b(49B), s=392b(49B)
  '{404, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00fb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 352'h208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 384'h6ac17d71260c79f81a7566124738cb3ee5d0aa690e73a98ae9e766f1336691e500cad51ba1302366c09cc06b8f7049e0, 384'h32ca965d6d7012ec187c7cab9544334d66c2a7658ddefa67e4ad40429815518ecc87b1492ddd57333bd2300b4660a835},  // lens: hash=384b(48B), x=392b(49B), y=352b(44B), r=384b(48B), s=384b(48B)
  '{405, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00fb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 352'h208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 392'h00e19a4646f0ed8a271fe86ba533f8be4fd81bbf4674716f668efa89a40cac51eec2a6cfbd92327d25efe91ca4ff712bc5, 384'h4a86b2e8e12378e633dec2691e3b1eed4e932cc48b28e45fa3d464cc0e948c02cc9decf2bb43b25937fcf37e9ad86ef0},  // lens: hash=384b(48B), x=392b(49B), y=352b(44B), r=392b(49B), s=384b(48B)
  '{406, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00fb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 392'h00ffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 384'h15aac6c0f435cb662d110db5cf686caee53c64fe2d6d600a83ebe505a0e6fc62dc5705160477c47528c8c903fa865b5d, 384'h7f94ddc01a603f9bec5d10c9f2c89fb23b3ffab6b2b68d0f04336d499085e32d22bf3ab67a49a74c743f72473172b59f},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=384b(48B), s=384b(48B)
  '{407, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00fb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 392'h00ffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 392'h0090b95a7d194b73498fba5afc95c1aea9be073162a9edc57c4d12f459f0a1730baf2f87d7d6624aea7b931ec53370fe47, 392'h00cbc1ef470e666010604c609384b872db7fa7b8a5a9f20fdefd656be2fcc75db53948102f7ab203ea1860a6a32af246a1},  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=392b(49B), s=392b(49B)
  '{408, 1'b1, 384'hb526d8394134b853bd071719bc99d42b669bc9252baa82dcafabc1f322a3841c57cc0c82f080fd331b1666112b27a329, 392'h00fb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 392'h00ffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 392'h00dd4391ce7557cbd005e3d5d727cd264399dcc3c6501e4547505b6d57b40bbf0a7fac794dcc8d4233159dd0aa40d4e0b9, 392'h00a77fa1374fd60aa91600912200fc83c6aa447f8171ecea72ae322df32dccd68951dc5caf6c50380e400e45bf5c0e626b}  // lens: hash=384b(48B), x=392b(49B), y=392b(49B), r=392b(49B), s=392b(49B)
};
`endif
