`ifndef WYCHERPROOF_SECP256K1_SHA3512_SV
`define WYCHERPROOF_SECP256K1_SHA3512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp256k1_sha3512;

localparam int TEST_VECTORS_SECP256K1_SHA3512_NUM = 322;

ecdsa_vector_secp256k1_sha3512 test_vectors_secp256k1_sha3512 [] = '{
  '{1, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 256'h59f100a7e4a774cf8f04577ebd9ab9ab2f09cfc5a6be10ffd0338524e6c26caa},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{2, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 256'ha60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{3, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{93, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 272'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe60000, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=272b(34B), s=264b(33B)
  '{94, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 280'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d4970000},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=280b(35B)
  '{98, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 272'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe60500, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=272b(34B), s=264b(33B)
  '{99, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 280'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d4970500},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=280b(35B)
  '{114, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 0, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=0b(0B), s=264b(33B)
  '{115, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=0b(0B)
  '{118, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7f68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{119, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h02a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{120, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32ab66, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{121, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d417},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{122, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 248'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32ab, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=248b(31B), s=264b(33B)
  '{123, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 248'h68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=248b(31B), s=264b(33B)
  '{124, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 256'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{125, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hff7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{126, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 272'hff00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=272b(34B)
  '{129, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{130, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{131, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h017d68757ac197624ae5c77dfa1b3bdda5c3a93710ad3a9c1137198b5a1f68ed27, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{132, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hff7d68757ac197624ae5c77dfa1b3bdda84e4b7d434ea95b99b774ce407efc6aa5, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{133, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h82978a853e689db51a388205e4c42258f705a5d6020e042a88b8d332b0cd541a, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{134, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0082978a853e689db51a388205e4c42257b1b482bcb156a466488b31bf8103955b, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{135, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hfe82978a853e689db51a388205e4c4225a3c56c8ef52c563eec8e674a5e09712d9, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{136, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h017d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{137, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0082978a853e689db51a388205e4c42258f705a5d6020e042a88b8d332b0cd541a, 264'h00a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{138, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h01a60eff581b588b3070fba881426546524653ea07b7d32f77af7137f4b9aa15d8},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{139, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 256'ha60eff581b588b3070fba88142654654d0f6303a5941ef002fcc7adb193d9356},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{140, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'hff59f100a7e4a774cf8f04577ebd9ab9ac745af2def77570c410612698168c2b69},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{141, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'hfe59f100a7e4a774cf8f04577ebd9ab9adb9ac15f8482cd088508ec80b4655ea28},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{142, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 264'h01a60eff581b588b3070fba881426546538ba50d21088a8f3bef9ed967e973d497},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{143, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d68757ac197624ae5c77dfa1b3bdda708fa5a29fdf1fbd577472ccd4f32abe6, 256'h59f100a7e4a774cf8f04577ebd9ab9ac745af2def77570c410612698168c2b69},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{144, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{148, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{149, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{150, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{151, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{154, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{158, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{159, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{160, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{161, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{164, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{168, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{169, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{170, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{171, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{174, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{175, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{176, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{177, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{178, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{179, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{180, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{181, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{184, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{185, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{186, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{187, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{188, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{189, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{190, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{191, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{194, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{195, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{196, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{197, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{198, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{199, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{200, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{201, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{204, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{205, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{206, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{207, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{208, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{209, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{210, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{211, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{214, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{215, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{216, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{217, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{218, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{219, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{220, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{221, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{230, 1'b1, 512'ha4efe24783e6e6cef1076318a92a899ce692e538073d95988da85c5ba8e97e3604babe2b714dfcd81aab90c522493c8a2683572245e680d13f802faa8f55ed4b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00dd1b7d09a7bd8218961034a39a87fecf5314f00c4d25eb58a07ac85e85eab516, 264'h00f5133b41774a185247720d2aa5d8826b6ec5af4c076936c8eaa52ed6cdf59408},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{231, 1'b1, 512'h0000000097ae34ada66084471ced074cb11f6012595501e4f88b5ab4526808fbaabfff3975c6cf53455cee950965a5b5b71310c8a1822cb5d15b513b43dc5720, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00904b2bb6e9de8f73243fa7ecc19a5a9fe034acad2b75b97c8cc84a79c5f35774, 264'h0081452342987040d43f50c72f2a5246430aa7559bee6c56663fd12029507a915f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{232, 1'b1, 512'h4a00000000d34b9c928306129f1a8059b199049f30ffd4d5b9747c848b197497634fb5190298af2f6a90d273164d68431c984e0fcd3a810ccd7b95b5e0dcd21f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b08122f027076f924cd1dc877c93659ecf942410772fba58881c9109311bca53, 256'h0287a0033df7c069fbfab7faefffddd7121908fdef76c04a1a402d599f04942e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{233, 1'b1, 512'hf25200000000600b35bfa47958845baa9428119e3a1641db59a3b72db0b47470dc44921ca1826d81bc2e78142986441cb6a6c15880383e1ed77282f966ad17de, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h48c044b94de8809898184e376a8a0903707679350e37ce290f858c8beef78c6d, 256'h6ccd83394e8abf4df2a40afb001ca4284d913d6b9caf6ef225d66bdddf9eb45d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{234, 1'b1, 512'h9e93cb0000000075ad177fa53827e2d0b2d93ab1e6b099c341864034009c13d5ae494352e6106d44bfde1e40f82fe0bc542154fd54365234bd13e0a0e4cbbf31, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h05535fc39278260eb2b8cfba00226cb3155d75c0cf6b418ac56df63b7c0b1e9b, 256'h31aebd43e848874347b38ad64ef172fa315fda09645c8752c0e010152e43418b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{235, 1'b1, 512'h6d22e20c000000000726c9469eebfd2e764c9b4750557869e51bef687b0b07862ad496e4c6a056d46f5d244f5f10ad0005ded39047ab8247ec969c4e42ec2219, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h78957c4f5a000af05fc477cc813cc6dcd9445438215b1c493780b6ccbd39a965, 256'h67023127ccde416b92cb3a7560436950ab643bbf08383ec9f4f6862cdb302095},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{236, 1'b1, 512'h5a5af3265a0000000025640fd363bfd88cc171f1966b1906138185d763f0ee7065ebd2a5813b79d02ca118763c60dcbda580f5ec322cdfb2c0a407e223f6b16d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ea1b7fd5ba10eeb70a456c149d494fa3757a209093c4dfcf03730d1cd54829e5, 256'h3cd204bb84656435e3656fa5e76edc4df3ee79615f7f1adfaf388a7eec4f8172},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{237, 1'b1, 512'h6c0f86f08b1e0000000069a0652407ab389f7f275bee385294bfc2a7a9119905f5ce4e1af41b3850d665c942f16914cf903717ff47c4e186c7fc97496a068b91, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c9611952ab603753d0601e0c97de91a6d2927d38afeb1b2b622ea384968cbbe8, 264'h00dc32c42ce627f286f7d14aa4b037588abfc202b916a7bf9051c3d0527c66dca4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{238, 1'b1, 512'h5ab9d448ee67ff00000000baa93e38832a2709f7238f9bceb67b53fea917f665de9153c44b7280e1a5674dee745f5350bb3f2259ea084b398cff74d33bded951, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h12c960e3fcfee173335123fe15cd7f8c8bc55f6f84a071e440b0e418cc9c0c2c, 256'h3f494246c0889b4213150ce77b6f5f2957476d3faf898135d56c145fd3af35ef},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{239, 1'b1, 512'ha1eaba175145939e000000007804c10bafa1416c6dc9d3311f844fe42868c6bdf283b946814df78822f198d26d886ed4713421a20dddcd82a21333d922eb39a2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00dc921912a76a225819d4956a7ff0660bcdf695bdf286288858ccd5a260012771, 256'h6bc5879138b207c3e4e692d4412c9a3fdff91ac58a669ec830b68b1cd562e556},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{240, 1'b1, 512'hb1fe8fe86f9994808c00000000f313a999ae7b5281bcacf933f05e4c8d526e761afa3141e9efefe959438620220c28bbad7047a6c1a98f95520baeb1d7af6278, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e31a34cb647ddc65b03f9bd05aa3e5e62a800c6fb56794843b606f1f08890524, 264'h00e7f2e4ff291bd309b0617478da0fdba92535376a69dc43061783b3ef928113ad},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{241, 1'b1, 512'hfa3ef856182ec646db7300000000241a0e98fb88ce661de43bfd86f1c929391ee9ce6c05612b1609d6b8466a9c4d0af24ccb440f463cd18addf4674adb2f94ea, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h47b825bdd67cb5d91f017d52ea77f59b1de1e05be48a469978fc88ca577dba2c, 256'h53ee369d5b89bf58b3c76218b7cecf12de68127152917c58ee155ee85dc664f2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{242, 1'b1, 512'hed19e69c6f4de76b35ce6c00000000ad94175b8ad5f1fb69995d7d87abd893772b81ff83fd6caa25d1fe69b0317ec4068cdddac49512e6bf12d9cd8ce9a951c7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0085b2d5faa65cd162e666df35beb535c797e7a2a20836d351ebcff798c343309b, 256'h196a837aabc19fa4522c5fac4c8e63e7cf3a5819c97fcec10e80f33e41f266a2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{243, 1'b1, 512'h2e2e984df4c5b45f7e337184000000000600f130d66940e8b4c0c1030e71fb8df7efce69100b9174baac3e7c474054e875f26cc182e925a17f55688964033e9b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00de538dcaf220334aca9fbc11d1576643662c66585e268bc0eb331608ad9523ed, 256'h1b1d32790d46c6925ab909408170839f83e6a03a7632ec8877a0c191fffbee79},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{244, 1'b1, 512'ha8f658c6632e4f474a6f1af1b9000000000048ac2a6121c8add714fb8cce854dbf1871b07a75008a42baa6cef01b4875eba4bc9327b41503cb36ac20f9354238, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b5d45e7fe1196bf5e076fd76742c1e12eefa7934de826d7395646c94a8013fbc, 264'h00f5475abab65d9ef64616fde95b3ca6b75fa864758950015441a4414acdd0c894},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{245, 1'b1, 512'he89af705f005a4e1c5983824150000000094795c26507ca965c1eaf5782dd829a5fb5464eae46688a19ca7fe5851291f76fcd7f7226131d74cb4dde6063215e8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d973f8f20c33772413f214d1b8709cceaad159c9211ccf337e7477da197d4953, 264'h008d4c39ee66532e2ceea2f0861ee02781ba0339eefb30bc06218f4a63fd86c11a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{246, 1'b1, 512'h9490ebaece67e31eca85b20871120000000077b2785e29958e0ab90faf8fcca953b142d51892ae5362246dc07a066ff6a4c9fed90a79fb59abdb7c8a888a9652, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c487ab066b8bdac12b5c728586a61e42d0a1bea16fb544d3bd56fede77bb3db9, 264'h00d27022a17957dc23bd760d0f00e93f10189c67d32a9ec5489514f140e49272d3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{247, 1'b1, 512'hdf22c290212fe9b66a9c65575e7be8000000002b9d4a3251cc7b64eeee3e76b7e65ac253a2e3d18658634eacb7494688a1616feaa0bf8a6cc0edbdeaa4533490, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f7777648b15af89af40cf9ea0a3c875aa0d9d736eca529af4eb6238f78a562d2, 256'h3b70d46e1439bc5d941bdae8507625971c1c64dcf4c51bcdb43b1ca3ae0373d4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{248, 1'b1, 512'hca6a7cd52432b20d8cc73c4e810dc325000000006ee638ed6bda85ccdf3b4606a300f2439910d382aa47f8e5839698e4bfa1756c5e93b3d6aee97edbc8ae7794, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7bb4646c887062a6c3e680b1491854c4b26a4728e5f2b2c1cc3087c780dab7b3, 256'h62900f55b885617f9b3c7ef34c67ecc37bf78e11a04cd6b9052eb80f9756559c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{249, 1'b1, 512'hd912418a7d72e83ab66eed185bd627c70b00000000a88db442365b3ec21269abd09b4b2e040304518850835236add11fecca5a2c529f8bc4c06174a03b997830, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4a96ed67d0950d97a8675c302f6102215ce0ec837ff53fbf06b57b010526b574, 264'h008deb5f7a7c8cbeff01c3443700b8da129088771c8c2bf4ceca2a5fa81138a534},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{250, 1'b1, 512'hd8cdcf759b329e28b173d8582d7a91bb2d12000000001faab0678de44c1caaf5247d111c9e465596a89073d5492cadb0bc766620952c817f31a391f32fb27346, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d9c3938a4b91d0660f6ddae8540a7bbeae2b0d717bde1f33e690428019747193, 264'h009b022d6547abf9bef980bf8fd67c366e234eff3aebee58a7ee56d335df807a29},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{251, 1'b1, 512'h91f07f1a3d4b600628f1754ae5ec28d43554a40000000051e8c4594c5a2e68bf2f497bfbc7e703e1b18398a0b5515a38d60284b1a2dfad8c9132a7b9a98db6eb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f855a2d237016b1e0ec307672a793668b611d2b6d4e5acfe2b2088aadd6296a7, 256'h13c60acb5e6fa51f03ee8cbe3a220f3ac1ce527daee05e9d7430343030dea7e7},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{252, 1'b1, 512'hc6208a5a5c6b71a957477d8c39b01e072a65ac1b000000005c6ec3ddb8ce20911bba1864112d3407082c700820f8676037efb40be95619c9f686163a4d0cdc5e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b8ddb1ed6e80056fb9cea2590b1b63cfd1e8098c27547ec8c6cacd78e6ebfddb, 256'h7514ac6644955744946fcb5617f8b067850a3ecf829d821f18435a5e11a4a58b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{253, 1'b1, 512'h7da7793b2bed3ce23ef7f1c04376791fa03f741f650000000008744fe10ac37fab4edf76492a339fe79e56ef75aee6c3169a0a61e3cb27e74666a4fe4184526c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e903b7ead454ff8de871fdf67b6bae4ddc88254c35b333a98ba3a2f6562678a5, 264'h00f713e10293aec60e63c2a79b189129e54919a74cda6a204a2727c13bb63a25ba},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{254, 1'b1, 512'h48cd33f55583315ab2131d5db1f9cfcb0590b13a266700000000c9bd5d6fbcdf457e3bffd7b4875145a47be68b99a201b93b8685e80d61ce692a913be1183569, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h615208d06b392c418fba55c752fef7b9ab8ed47d98f40776d86ff4bfa3e95464, 264'h00f403d5984d446acb203eba58a5468372267f9004f263aaa1eaa208652297db5b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{255, 1'b1, 512'h1acaa001f6ed1b1a5b0bbde85513fe0b7aed266bd9da3100000000dc1113ab87ae3bf815157a1926b7bc3f659934702113570c26bf1bcdf1c8492f79614e844c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0eb65a5bc338cd920a174648dd84ed5443f37417d8d730ceab0dd3fb9a2046f3, 264'h00c7a86d7e09f5e142fc6d45a136b4581e081f66a26fe0255f012b812d7cf90189},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{256, 1'b1, 512'hc6244ad67598a847488d31d513fc9dbd21d96307c296a4170000000012f527d2192eacdb6045c48c250e317b7fc62ea79321783ae0f400ea4a60b48c2a2fc495, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h226464501f1ccc32f1e1482fff4624f4949343c79a820d4b9df637b493ab5b23, 256'h4eb47d0fd14db448cedd611e1dae972bdf27ce0fcfc19d9ec5bda9683081598d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{257, 1'b1, 512'h90f9b7739bb1699b90bfdf7cef079649e3f08242a08d05026100000000d3a4568eccd5ef4d94de4885986b68670617f552b9cb2a6eed337392b49ad4d04a9dad, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00bc0d706b5fdf102805cf83f66ce17a97aebd5e3b6e7d5c008cd51164750af108, 256'h651388d190da29748df343dc61e23c248c753013a5688652ca43d222edd1bfb4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{258, 1'b1, 512'ha7ee711aed6f375a8a15680f30deb6946501624b70b47c79d5a500000000ee6f7f0f2b69cde1a389e3abe86e51efe844c8e4ee7c3b2a15925d8c9b8b296ccc53, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h39a1d9927356d6849b7e96cd34a5828bad112687198637e7b84900ed92fad0b7, 264'h009b5c753e2e10619e1993b8d8171a7aa4c4813a8721aca1f79bef06c0fa858462},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{259, 1'b1, 512'h9583a32b620d5614a1c36e06ee45750fd69ef561faeecded2ff5b4000000007bb68b2b419fd574ffe1760fa0203fb1718c4e5d8a798563fdd98439f37a56dab7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d57adda8926a6b75a5c994a0b8abc75534e68bd79b02b8eaeb1a7add4c5c4232, 256'h3b349431e37740c60f92c55dcc8a9f55e70e27b9f73d82e37d728ba7266cddf6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{260, 1'b1, 512'hb6e404060dcf7182366941e77a0f0b43737232bbf9f73865863c271800000000a4ea51e31a92eede7497562eb5eff19b08310fdcd46cf3c22e069110aedc21a2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d5b4c29599e97085686534f843d71d25f22b96d89c70b4030abcbe6abd73559, 256'h28797ed87120c4bf50e37b0704d2d3b4e0b1b98c27e618eb99568b08123a1be9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{261, 1'b1, 512'h57003aeb6ad8b84b54cdddb9243c65d8fd07ad1ffdd35f11c319f06394000000000aa9393490e8dcaf1c1e53ab5a7b2dfc0bd1dff4d0fc1e0c9dd5cbb035748e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0db6c547a1e7bbb715b48b7974104b6d7618f1dfed77019daa29bd59b273c087, 256'h57f054587cdd5628772c14dde0a77dc5c1bad06828410c5c63b9c1b35fe04410},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{262, 1'b1, 512'hb47f61cf42394fa1c4c8cea80b83e366e30a938140f793851af87bd3782900000000d7a39fae605c98c96e0a5b0e8a58e47c3b50d4905171c884a64239fdd901, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h094a1e172012d9367852f228f49c382bbdf19a6b354b8511807e585cd46e907f, 256'h0e50740da30419a987ccd56746b8737aa74a1292892eef99a34025aebb6dd209},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{263, 1'b1, 512'hdfe80a6b887fa09cbdc8bb94300a4ad38f0380331a18c0a0b62708e590dd3800000000d364091041bb72f35391e792802f5c23fd676d0775e56ac2e41880d92d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h73a5445895e0796686dc28c3e4cd5bc1f85368b3264b455d470a7cbeb7592d91, 264'h008a9ffabf9f65921734934d65053a00bfa3c353ac81cc9b6f60271635026cd0e1},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{264, 1'b1, 512'h16d0d407630fbd8dd9af18abdbdb902051c86b156254ecde6a5f0a5a1510f99400000000c202a44b1c172e1436f2252d80f9ab44794b22086f877c3bd4aa5fb3, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0630f2c6277e9e0414b7e8da64311850b6f3912193970fd6e2f4df79df720c7c, 256'h6ccdaf47a44ee1043b76ef62b3de3aee876c26f4efe492cb3649423e599753d0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{265, 1'b1, 512'h519e4709f22b7ec44e321f4d403bdde7f532392786df003ecda243880f79f899f7000000000e3e6d749c0a602d959e0fd13a8a491554d233b9dcce6cac4ff3fa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1e1b75a3495bb5ceb2adb84b80f117672b79c5bc71e953d1a274b11dc4238729, 264'h00dcf48d930d89c0d301e97f9083487e63cb39127310b0f5e3c8769e98e5b2605d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{266, 1'b1, 512'h00ac9e66bf4db08b47a08e0b34e95e7ec2da8a82091479dabd2d57199b450dda70f8000000005b979f8077a5a74eaafe42ec70504f2bf8cd07aa23ef52c0321d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb92e1a80ad7f440d8a2e9d88ac765c5cbf724bd367f414c9d91cc1904afe497, 256'h74fe0ec7cc0122eea4e63c4d16c89edf6a57823178c3747b01e7aff3df710007},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{267, 1'b1, 512'h2cd7eb20ee13fc351891dc4acccbc978161cc1b1e0cb95127485ff132176a972377cdb00000000add5eee3b407ef394da0255f21b9b8ca144d7e76fb075c6bc1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7c99e1ae6941f4bcf54ea65491cafca180eee1605a2ed908c476ee67cbdd7373, 256'h1f94f03ed47cc9674abb294cfe7e7b10ad67101b8cb245a8b5fb883a21a06dd9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{268, 1'b1, 512'hca402f2de7f990c5e1deee30d418810cd3a8707888fa5d54d3a5a0b3bab20144dbf37f52000000002a1f22f563f07cc9d066dfa8881777cdaf8a1ae4d43d6341, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h29bd14a9dafbe562e0c4c0d4aecb6491bbd37f707133f78fc5cb3313365377b7, 256'h2ea1d86246d8edad31132f3dbe642cac488690849bdd7438d5c626cf8c973970},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{269, 1'b1, 512'h4386a89b56a955feed663fb88786a1c3916e8c65775648439638f2278c7d32c6d67f942e7d00000000d3a5ae2110db187684130f7aed62cb05159f8bb6eb1b26, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00cf7219dcc18e22bd487b6f59c6494f637c5f0ccb18192e9e60178621220b49fc, 264'h00a05d5abbe25a610c8e3615cf7d01c69563ddbfe76d7235fda45f046af03e50ff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{270, 1'b1, 512'h9a76ece71e15ffca113598c14654fea437156151bf5c8d47e15a6279ff965eedbe79fd4437f300000000148cc8ba720cd12a6cafa72448ec2cd6ad2852b2f703, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1589de61cd315ba0bf7f0e577f00589d28f72131f4c7af41c6bb31ae8ba271da, 256'h2ff82a9a1f52901c4c6f8b8a41c0f6e760f160da266d788da5bdc945084dff8d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{271, 1'b1, 512'h24abce8b935764d6a61bf597db6c773145d5992485866070fe22cd0f6f871d53e72f6abbcac6ee00000000840dc44c1955185bfcf393a1786b04625904f03e85, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00a8c59942907039886bc374c17ff452b604385c3537b9b6c6113c1b19d72e68a9, 264'h00d376bc866cc82d78ca17b461edf16faea44e577659b1fef02cec0f41bd2e747c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{272, 1'b1, 512'h3fa9e7c5fd635a7b587b56e19e8921e7cdc6d8f6b1ff03b579b907ccc2dba540c1782d5c35e3aeeb00000000a610ad03b540240313bbf54453b27d3794341d59, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0099cc652412dcdfc574b6fc2525615e6711caaf7d558cc781a3a11cf371f40f71, 264'h00866dd4ab6b58b5d6379f0b431f9a251399defd5516bf6bb5495511e05b24f801},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{273, 1'b1, 512'h4025a46ad55fab109832d892d397d6e50c9c0aaf7136c275c259a6a61333a7e139b394a288148e32c200000000a3d26314f0694c5db5058ee34dfdd8fc2af9f2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b47cad5c88161e29620957061e24cdf46f3fff97c266b1635fcf2e9cb4d92879, 256'h13549f3b1b639eeb33f40cb338ecd089b9094d9625b76734f3803e9d40a1eb26},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{274, 1'b1, 512'h1e2fbff1179de8374cc3b5f47b00ade36b6494b8941aa810476c8b40e3ad3d7f5f60d8ff0d13bdc7683d000000005b2a7c0d9bb60d8af2267c656e800069cee8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f4f3a043b5bdc56bd471876e2df15ea80ccb189b25486e6ab9007cffe121acfc, 256'h78e8e3b3589580dac1ce299a18f5704901104cd21205317608c330adc8d35272},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{275, 1'b1, 512'h1efc0d2c8682584f2504efc8fb5fd2848583ab11c97a1ad1d23db89d7d853316fd159eb4e2cee6ee4f2eae000000003ec9bbec801c26e55e61dbd6364bed8027, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5df45e90f9413908b47f7cbb05d6c43a81eb62375ab961d2b065c6118023c018, 264'h00d720a2a23c34ece3acc1a516070bde6bfcad28fd89c482d72b69d8113b1903f6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{276, 1'b1, 512'he68fbb72e90ec509836476f39f26d3f65c5deffafd5b86448457438ee0c621fc8f97e83c77ecd131ff1e33e6000000007c2a942574c7da923726d5304e0de79f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h780bb93f52d53752a9a877dab0578c7702d1ea889960e1682e84f82740b1be5d, 256'h08e366ffe8f72d041426aee57aeffce7822b209c34b28255a5de67190870ce42},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{277, 1'b1, 512'h90bc23f7e48f29ee5cf5bda8b42a6a8aed3cb6018636758be3051cee87758ed5998aad924516e34c49319b58cf00000000b7f0c29548e1c1244f0caff38b285b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f743a77c86dce094cc265a87b2e053c8cc773370851dbc7ba1a52c58df24d554, 256'h2516e4614dd7ccd36a23cbbb1b58c29f900d4da2113e7b9ac956bf8879907680},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{278, 1'b1, 512'h1c0e382d29f7ce824206c57f19794f9e8abe01e6af45a57dc9c01184c7b956aba27c6536c48c0951e2540bf566ac000000006db962ed4d45bf0d0c1c6c806b4c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0b77b2ab21a5c92cb0e3f2f5b8594edcc0dd6c70dbeea9d9d363a3718c64dfb4, 264'h0091c2d6515ff6f2977fd0a150cb04c600102f0ae07a9061993244783e62f2337a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{279, 1'b1, 512'h92cc3187d3326341d51f43165add210d496557c7a27669692c21c2912bc85d13d22a15ce9f2dc8052f89cdb3444fb400000000da250c8d1d81c198686e0c62d4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h41f0a220d11a014dfe43f89ab647abea430cf5a9703088f28c1222abb77e8857, 264'h00f811c584c10a25fba6216113698e5a2dc52d8ea340d92ce7a11d356f6d5a1382},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{280, 1'b1, 512'h0ec91d81506646053327c352b11803f36a38ba32d940cdec35246744477eb4c423fd81dfe4e728bea623290a65646d9200000000f68a3961185e3a1eb3a74496, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ed707e3cac8bd56a4f0a3118558e8402dd477be7dcaa1a7ff448b0bcbfc0fac1, 256'h3d9933e01d7e9439059973fa499c37b896213b04346bb292f867ff3a58c3d07a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{281, 1'b1, 512'h290ba1c9dd4ce7537613a8092317a721e35cf33f17d8c82bc20a765683871857d7a7f0f72e659928158b11760b339f16fa0000000065c91469026a04f6e368f6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h008035d10dfd533e01718fa9d0a1773e55b424770415e570aef766ea2cbe577c27, 264'h00815b0f14d6f7f4ca45191428d98c9b414871ffecdac3d0717d285a473e5ddb06},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{282, 1'b1, 512'he9caa5454fd145db00275838ae34244a94ee61a025a174247c1b8056e6959c7f851f3038bc773457c88404c0dd497580644500000000719f683608f5718616e5, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fbc3576a648ebd633152fc896ae6b4827c55824fb0c96fdd217fb2cfe3bbe636, 256'h0b37a95b15589663db322e1f089aa8132965ed6490362d243ef749c6094527f2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{283, 1'b1, 512'h1827524c50d2a178cca81cdd33a0be182f764450e04af569ce80811e55ddf11bf9b04675631ccc24d816b26e407df93f288bae0000000040fb10fffd72f8f6b7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00de08cc84004d3fb30521b8e0ade66b6d52734ccd182cace8a34ba0e390fea893, 256'h2c1e3deb79d16117ed84c8982276d43709c5963d57bd2b10a530ebf161da1a3d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{284, 1'b1, 512'ha5186acc06258c75ebd6c4985b00ae514a23405ece5e1c0a51122b5727c5b17a8adfca46c2479895b4121c304b5b2785c72c06a000000000ded1a008316d23dd, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4eef795dc7b17efde95dc52062e3b60ab360d37704800fc915785e7739b834d9, 264'h00c68356eacc3509bf4d2b62412b2472f22383d18fa8851527294b1fad194c7bcf},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{285, 1'b1, 512'haec77ef7d501e59ceb458f4b03194d730583d8282b6bb01ce0b0417143ca15c2059e8290afa26d6c1e38502d0b895bb4cb182dd4cb0000000097ca7caccc470f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00cb845b9fcfa07e88e9011f0311cae9f3f740516e7d16d9819b7d0f6fc764dac7, 256'h3d7f3ba5173e130937b02bb7b8da25c506ace6182b8f9ae4ed891f7d216c0378},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{286, 1'b1, 512'hfac59bb2cb17756c53956cbb809fb1dcf8f30340a8b21f7a25a1e6b500284c29820250c5c8492ecb2f1c5906b55dfabfb8c47b418d50000000000efa79a0e20a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d19ff3efc71258f747e74d76f091107b1fa47c87c638720b55178c0655dcbcc, 264'h00b8a653e31931dbd2ffc4e957675c68c28719b8118ec3ed3778c57ce3eff1613f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{287, 1'b1, 512'he1942b44674c9c247d1f5857111e24baa87afe02ae74ac9d1ac122c10ced967b6243fd3055a4de1d50b98e24831c9f613d767a3060f7f600000000e5461279bb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h10d465e03829dad77e8246ad11caf8c6aa8aa918c2bef5a9a9e601c5a919f68f, 264'h00f365a7a7540dcb642de90e6d6ccf0c74094a8005deaed4062e394e1cf2bcd8fb},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{288, 1'b1, 512'h9ea149f211e7bd1f624b20fd50fd2c474d627b16250fb6281c6bf57af0b868f48101c656162b5e1415c87cbb7a685fd752937f97cf58a424000000009deec0f0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h674330ea5a5d45d71fca1f3ba031494dee9a8623e0d9e9adbb2822794acb4f12, 264'h00ae4d3830157c820bc23fa792188b94bb559c3a6212768d7ac59dcf36f74402f6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{289, 1'b1, 512'he2d392cec1344167d947974fed90e637c5f80aba4fb00ba57dedea9f7ffd1b0404437d90e50f742cad5ed8b82bd136d13319934da1f04f50950000000059c93d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00a632c676f667669bda1b0ecf5f33fa67aaaf8aee46bc9e9f2bd5bd10c36cbb95, 264'h00a99352cacd6bd42b78a93908008c23eec2d36e5e4fd0aa349d5634fc543199c5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{290, 1'b1, 512'h40195fbc1bc4b600980e2c2b763857780d875bf68fa15558b038d9333a6c76f3aa4687e0325e29c3945bb8ac11ce675dff92bd5dcf0efe1264e900000000cdc7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0c9d2e8935f855e69dccd877d95248303e1b6daf8f61da500150185f5565fa97, 264'h00e4ce328f00e218aa13d496d85b73b5b891cf0b7c66ebefe5e6b92b1da7f837a9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{291, 1'b1, 512'hafc1cfa16e5549a03769a98e0a323b3ce3d8e3f316cd9f1007e4366b81a3affe3acb663d6a5d6a6857c736ce28eb85c432aad5ea98a80abb0b973c00000000b6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4748c00f44a6b3a8726f604d7b933303d98cd458b850ff2d7cb90c11d5950ac7, 256'h766df7aa4c8b3f8b03b0eb8aec653fb70eab7433a84e7ef2d57f368a051b704d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{292, 1'b1, 512'he47ec71fc0cae21e08260f64fa9dc1a4c99ce92048144beeaf932a124c0f87a8b0db214e5424891f30a4cc0311efbb2d49807cc31733db9bd80f912800000000, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4e4fee37b0b93d7d6dbee89b47dab0c065186ee81caf2227bb26e85149bbf9ef, 256'h3eb83850edda9a1b1011118feccd03e47b3e1ec815837bb7f8867288ad8df831},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{293, 1'b1, 512'hffffffff149aabbf287a78cde6477453f7f9c2310cd2d58ece43bb07019c69c965ca25e8df7696c97ee4ecd4966f7577eb41a60745d031a94f5856e1a5f95aa5, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009e8520c5e8296935fe93da2dad55963b9f1f88187f76810fff53c0a6e95b0c07, 264'h00d185de4f682a97d28fc3067d56a3d24f743f32d47a6f390068b2ceb71678fadf},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{294, 1'b1, 512'hd5ffffffffa5bd8691d54adc06abeae7d4857cd52aa3ebae84fb391361d804a381d15d6fabbedebceef14c94b5bbcf1560bc8b97cd4c4accead9b453f6d27746, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3cacb67364a3fc1a379557f7e6f5d0f501977fd4822666956c9356146b7d922f, 256'h686e27be6217045a5010c88003dd3956a864798c8ae687714fc8b7277f7b520f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{295, 1'b1, 512'h9481ffffffff6e35dfab283e61e8f9a49de1cda44cdf1e2680292ded627b16d9b566ac057cef4c3380ee126c020a6ae86ded132faef613440c54185ed5986dcd, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5df702c77d4638a4302d21a9fdd70bbe31a4a4a79c7d531d4f4c8283970f664a, 264'h00f72d799abce3cd22985c5cfc68f7afc8f96f4e7dce8485ed5c595edc1e1f1d4b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{296, 1'b1, 512'h2d8fbaffffffffb42e8498ddf2697ff4a2223fac0c486f05f57374d84dab9e8d13f52f6c898c8a7a74f2d48bee3cc16265e12a6dca3bee77c0ff0ee5e9af7e49, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h243a857dfd167b938492c421bd657659d101944736fa79b903cf91ec1c49e8e3, 264'h00bab3f04f130d737993ec8f45503376abe816c2b8e5ab3decb0dbca4f5e181d08},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{297, 1'b1, 512'hae17b907ffffffff72c833830a0827c91ae711b1704754016d3b0ef4c8367a7e93d4ba6f63e6bb8d572c24bfdc55da0d39f5fc8def9b04723ae25c1b82a3ed86, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h67a7996b7680e958480ac2f97084f2055194b38e0ecf82246dc87918ee1954a8, 264'h00de187dfbeefce383dcea1a7fd71362385d09c6d25aacdfa34ea270a91ec97cf5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{298, 1'b1, 512'ha55ecf9029ffffffff0b0266df6f2fc70941d6389583046c5649a1740aae64600c31269408a3fe8dc0975b57d60cc95053b7d311b677bda6e8a0d6792e328bb8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ab6cf003aa7865cf8010ea01944fa0d2f825ac6a997a427f8a4e791e797ac6f6, 256'h28a7a6c80582ba8f888d2008fbd696799561e92d9a51922cc602aec2135f08aa},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{299, 1'b1, 512'h37837a8407b6fffffffffac5686980dc2ad1a556be4d1fcf5dc000a18139c2322fb6d35995be1b96f942fa8bcb31b6d4c0efcdb2febaad183b00f4967c63c04c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009f9f0be992fdd3e069167599dc55e331c9f189d2c230ae15d1b5b441d3843c74, 264'h00f8e5b4ed8ead0352e032f79b5f0475f0975e3738d784d895e9e4002b26762b79},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{300, 1'b1, 512'h148ae8a9d1f212ffffffff9007e49461386bac4123a9f847a6901d8d1508c822348ae29c100f38e169470e9a05b8cd6c780a06d49e062785dbdf1fd4cb89afbb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h373b8587777d2b4ff461fddf521abd8fc5d3a1caca847f4a5461dab6ba242d83, 256'h51a98da2628724018dff804c26a9671f7df3e24490392a2d1a91fdc7f50deab2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{301, 1'b1, 512'hc17991fc38743c0bffffffff12be8c0818873e8d65ea350547aa4cdc067cd0a4c21e1d9387ca3c60306f95160cc1f85a08ebdd4f3107b359483b719f5b9a18ab, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0090a6286a271d8ffa72ddb55e8c924793e03b2af73ce10f2deae857961cb07070, 256'h28df2b6379501110c12ac167189f9ea8873e1d62ffc76e6ada83f2cf412ea5d3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{302, 1'b1, 512'h45477dd24fb261b2dcffffffff376705fc972d1fc0eebc57960e96dbf0315340601ad9582193434f8cf1ff955cfa9a803a99d9465ab1d11337155273e65b2735, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h107434a824ec05568d52219ab3e847046f01493f1db57a82fabe754555838292, 264'h00d1c2f7c1ecb5afbc9b0e63e20fcf34cfc16bb260b0748343eb86c44012449b8f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{303, 1'b1, 512'he4d30dcc9e0b433fac32ffffffff83bb0169390c4443bfa7b7bc8a7c4421fb94a64d266b35ee622ee92a194a9c369a1bdd0961e4047a4fc3ed632b51f01547c1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4b737fb724c97348fb67a994e88816b1091951b77234f1904717ec7ef1aa951d, 264'h00ff722b669bd4342e6b856232b5a5c03d2cf16f09b3d3842d0a87fc19d910acd4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{304, 1'b1, 512'h8f46b06e493783b6d3209bffffffff5f263101ceb63bd0313945c63e59a123011230ea2a874c147574859882f49e6fdc842cbd97843daff440629f6a58573ee8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00abe804f6c76fa3f1470c0f244a7ed96807ddffff4031926cfad9a2c9f73ed773, 264'h00e48352653ccc46f5f5a76d7eb3997dfd412001fb1692312788f7c297ef792fa7},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{305, 1'b1, 512'h34de554e38945bbfefa7cde3ffffffff7b63c616e7853caa71db174d8c61626ec0c2d1fc20cbd176f51bd580fb3d6dbee8b1319ce824b44fd820e94589a562ad, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7d55a5da3201de5343703ff8ee363b7ddbcb3d786afca8f157b25e7c90d09de8, 256'h3dfcb55acd7def4218abd3f989e901f824cc2d4ed3a37b8794117975103ff004},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{306, 1'b1, 512'hc80ad608a993f311fc5d85b14cffffffff76d81aa75f097430416ac8d6d4e8f80858d995030cfd10467787a708fb59252ba27fd5cb768e2b3cf03a351aec1402, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h25d2c88f0b79f2289f92d3ecb6de119fab764fb43ab5286391f9a282c82ac198, 256'h105f44fa27afe4dc9800e6a16528314de01b17737e9741862f93ed0cc33b30f3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{307, 1'b1, 512'he9f4410a9857187394e0dbde1bc5ffffffff22ae4f317b16e8c82ca5e8ed1488b15705fcee61951d122b9603a8b3744eb429a850db99537b15bdee559ceb17b4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d725c2731a6db8d623027a926a665e9dba0f95e90a5fe6807a84b200111f04ec, 256'h346140bffb84731f0f1cf857193dea25a2f721463dc3b85a8e72c73ff72bda94},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{308, 1'b1, 512'hdbab4c37e253fc1deaa9e71c035737ffffffff6e927ee1da438de0d1d5152cd6d0549d2b8172bfeb94749da7ff020aa760407bc5e12a5a099a45a301588b62c4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4fa9704d3eaa5760da0b97abc0de1f872840e58bfdb1a8f9d8be3f96f950ca7d, 256'h6ae15b572c7d1a49c99e1aa54de5fb2bbe055d45686770f579c08ee79924ede9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{309, 1'b1, 512'h2ad0f69e7f2e5efe8116b4b576a322e8ffffffffd986d354530161e2776001b50987f4eaccd1eaabb1c1d4d6c94e4f7460ebae1ff8cbf4a1df1cbf4a3e01348b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h343353c8be35ca222a38771b19ff3550abe41b91f2ffdea9c9f4887d70b02782, 264'h00c285e3761c6645b3db4ff99a7ac40803286f28475ba28b9cd55cacdefb330984},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{310, 1'b1, 512'h69e08e9fa0546aec130be51f245d0daeddffffffffd8d24508cbc6106330bb7e4453fa88ddeeb7a8b80db338a7f66e078ffe0ee91d6b432c2d52b5a0a15f847a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h529b121d5b3cccb426189d7343d571adf05cfaee843669da6722f728c192bb82, 264'h0086490a7686215fb29b18a166bc22c1b8a982fd7d57ab593318adf8355684b45f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{311, 1'b1, 512'h21e7350eaa2b2a36fa211d7c6b144fc87b5cffffffff9c3a4d277dd4c34a428a3b35dc4d8c1840740df3876a387e6ae3c97b0a40325ae41007bb1de4338ded6d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ff65707177bb9aa135c5fd774bf72eb3058e80afc7d8bdea8f7fd18040ea9959, 256'h0d4ed13f9e01bab8aaaa40d7f5c923a78470888375b4690e1164a83fdf136201},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{312, 1'b1, 512'hffde6b2d174d86702f3a46946c7167cabd18feffffffff2df58cb555aad0b0df043b0c01b91bf2ee4827aac1d987f3174e1fce7921c831a0b0aeab1ad1156fed, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h471ebfcc45de07bd4118f94b0284f0c5848dd93149a217b56b49e20baf583ced, 264'h00ad498b79d6151bf64e003f502fca8fb7b05b2106a96ca1b977ee002c73bc721b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{313, 1'b1, 512'h55260440dd65e8c48db54c801af143d639f08a95ffffffff9f03419e88a5145c37a3193cc07c160404a9b7d489aa324965d89fc40fab65a71fae34c56afa395b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1e279add50ce6148dd4a3d311bad896745a169364ef68b94e6360fc48e949b9f, 256'h7230fbe4007fb7d6a4274c396081f37a1c9b2559b526db1efe435ead15e4b74e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{314, 1'b1, 512'h16438d031fffee5b56365cb1a8f4bc19eb046a111dffffffffc16998d3235c27ddbfe7f1e45105d70ecb963cf511b0e09daa505bc426260466ec6528fd48b88f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h52dfbabbcb99651021c025a308530b9cd04732f43463bbc51160cd542d9028df, 256'h0ebef4f6870bce1ca302e7120560e5170067c0fb3dc8668448b89dd4821b53fb},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{315, 1'b1, 512'hc0635b12b9164d0a9480ba133839afb60f79f6e7fa22fffffffff18d9363b5c503a5ae2f4cea06d8c5333965149a2cd0ed0491d1f9c8cfbf12fce9914dc22f30, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00dabd19aeb87fd56119a3354c468f4429fc14421c54e8be9e9b927941579ae55e, 264'h00b10a7396c973e052af2944d37247e9016682d4da7cab2d5428618ce120a21056},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{316, 1'b1, 512'had86d31823a92384efee57d7fc747fc6347312c57d7e61ffffffffbad8263d3a80dcea096adc61333c39ceb1a06bc016fba8beaac8adc0692127ebdaf8bb65df, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2b9950c4005dea8e603ffe0fd9b3f66b7c0f07509e50913bb825ef7ddf2e6e77, 256'h62c9fcdf79026f60f830e7cae4af814db2cb58b5a948562772da130613bbef94},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{317, 1'b1, 512'h155ee257be62746434e431f20477a5a614b621ca050d7f78ffffffff517e6eeec93db0df6b6358b1f45efcb67e7b201fe4b0f7ef4fe49aed869621bb74d2604a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h09d881e300448b9eac33c67f10c061c2c985c415a414d09c891847e3eec88598, 264'h00e75455a508493506f8746074f8bb3698d4362f98a9daa20fa916f6c4023764ae},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{318, 1'b1, 512'hde8b1dea4af73e03d31712528653ece2fa048092693f2106acffffffffc4fbe785cc6cb125a5ca069dadd2dd809bc3c6246bc299c2bd84aaaef1085a561dd79a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2db5a6d9b16c61c888a5de064f621e45227ab63efba61ef210fe4ef81c93e00f, 256'h04b8e57a7373b3642e58db0cc652d6da541d6d25c7b32c1ed2b408c9e3c39719},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{319, 1'b1, 512'h372064a97724ffe3dec873aaa5c4e830fcd9ac84f1c4edb9a372ffffffff621efd798449ba3d7c009467fccb63c6e9a825df2926734122b80e8fc9a6c956351e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7bd46dbe132d95aff854bebf1c0dd1e90303328fd84d381e93217723d1a4bc18, 264'h00f795a0c68d6c318c038dc37bd22d36bce8083096637e8912c3d01cbabd3feec7},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{320, 1'b1, 512'h0a55bcbb94c925c397b334ec37bd5216789d87fc6589738cdccee4ffffffffbca7bb2e94ddb13839ef8da502b39ac80f25abca143e0add021592ea7a36ce83ff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0ca03beb6d348d3d36d2e9f6773e5882ded66fe6026c9c27b847e34523c77c2c, 264'h008770b6f0b6aa7c982e84235f1840a6172386a41ae75fd9affac7916cbd19f8c3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{321, 1'b1, 512'hef503ce85b5b48ef35abff5d47345a71aa715f5e8e1568c9721a78ffffffffffe6124c567f2fb5b5f476271da455e079b655dc8c9506b65d9e3c60892984e8ba, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3f1a74c1dab6bfc319da38cde7a812695b530c60b36d2ae3fa11a7206b2031d5, 264'h00f07f8eb5825b2d5642443185d6afd2264e98996dc392519f812883dbe0e247fc},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{322, 1'b1, 512'h5f3afd4f98713d775d93b166838053fa503faf72cf3c00b3c57e0fe3ffffffff7b74af7667db987c9c205466e00679714af8467254f2e441ccbf1bdb9daad40a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1ae1c3ec96f8591a3a235de7c6f739201104381eebeab5fb5ee523f577b6c7fa, 256'h07ac1a9348fc8946964fbef0af11dc8b2da6feb3eee8cf475c4926ca9cd571a3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{323, 1'b1, 512'h9e670958749c5bbc0cacb1ee6c38e71eede821d75d84cc2fe1335af9f6ffffffff4e9613cec31f535c4c7bdab269d70a8d4b3bdffa3065d91435a4237cae96da, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c6ef5423c69541caa3bb8f361f4fa9caeca30fb329a0da806ea956270e0a9928, 264'h00c045de5205eb8bc861bc159522b41c0d66e62fac0f58730861000cdf9e27bd96},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{324, 1'b1, 512'h1e77a725c36046bc3bd6ca38747586093510952c0a3390d86b508479c0d6ffffffff25680ce9cd685ebae3cafde6315263f7cf4ea6117ccf870d42189ba3abb8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3097d229239b4085e3fb3188106d5da53456752976d2c4ba82dcff6ab96d1909, 256'h56f60ab76d33bc94ebae3042a1d56a731429f1bed162bf3ef7269d912aaeea71},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{325, 1'b1, 512'h59f9626626a34d5491d567d0315894fb702c1d7a2ec677a2b595a772b20d8effffffff20557e965f33f606242a59aea4cd565aecb931664e51fee93a92ccaab6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6c9ecb8dd5b8badd49ea1b26ae3ae2af7236cbe1c626aa6b27029ef1d6d05901, 256'h06c9bf356441f84215b006c721a00697cede6941a18fbc0f9c5b3c267eeaa371},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{326, 1'b1, 512'h001db8dc4aade36062b6ddb62bd342923f537cd35c957b47803909be234a3b58ffffffff0b537f24fbdbfbefce08b061b467fe60e7f86531ed3f54c6e29889dc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h43ae5619f91b711a61be076581f91d382c39fe53d500b136f81be639bea76add, 264'h00824594f08185479731ed095367c04def2ff196229c5b136b3835eb8bb819c56d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{327, 1'b1, 512'ha05bf269c6959e1000f754963c2ee746346fac0d57bb119d3cecfa3dfe702fef2cffffffffddcffafb72da48023b4eae3593eb7c3c2d758c1c6c5e4dc57d53bc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h13e8dc460a0d2af2305a6abfeac834737d4441576b194fe83147b7d7d1247479, 264'h00c590a7b7fd6de8c2d658aa2bde97de84505985e2979ab2a527658122cafaf61e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{328, 1'b1, 512'h9695a59c40d735b329f1f9c2ffd974ea8e66af6c65a1f7242e1eb02ea6721f9460ffffffffff9327209276e0633e07c96c9a2950a09411d1eabeda48ba90c8c3, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h27feb06a4c5bb046162467e523b4b62c2c8dabf26ded997eb0737d3eafd16c8a, 264'h009ce87c4cd6b93d1ec3b3c5d29fa415cf918edd24e0febd7b200d6c82c91e5f78},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{329, 1'b1, 512'h521abe64cfe7fa37251542760a99aba478c8b79a5eea4ba1fa859e6dd8bf23196e36ffffffff157c00247c6e0a683044034774f96f67cdea42afc9ebe8d78be0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009d76a05d5803a2da17dc2782ec469c8024b1d293a38c23ac4eeb3058595a24a7, 256'h226595b192ea8336faa44670fef5e808ff9911ccda85a1765c19ec44671b0505},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{330, 1'b1, 512'h56f7dac71cfda3cdc27537a7fef1026211918d8041d79637eee4bf44f6fda371a67755ffffffff1dbdc9ce7d24880544364cd8cd5925c287a256383c78631a0c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h791088736561f41932cd86f066cca6d63d4473aebb869bcc70c923ef80a7fd95, 256'h33402973e7a824602712a5abf7030bad2f183e6b4fa40c66399a14ae48e288e3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{331, 1'b1, 512'hba44f1aa7dbd00300b9d114936943eb2585a2ca6cd8f11fd68794b5adabdcfec1919ade7ffffffff099e11a571237729c09fc81d86398317874c3722999b1875, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h52685eef5f2168598c294870188c043dff0496638037170763ef5778b7b6fc1f, 256'h79a88d3e7b2c3a44be4b3b3305e4bad5fcfe07d179136f5ac926315ff9d4787a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{332, 1'b1, 512'h125406f9b34e4f63c0a2288bf6166292074a0fed2b2c47822bb885520f2db3e2c58186b926ffffffffee3b259d2c85d9ab10b9f10f7f3cab27a8f528b4a82ad8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5db883b5a3766a2a14ab26a25ec598f7bd1f97585fe0b55341e7da251a62ec1e, 264'h00bf63c66e992c91fde513abdbd59b4f9f542881cfdc2be3fbf3e772b97e505b3d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{333, 1'b1, 512'h46943ed052f77d2e9549dfb8b9a4c779959f7b0a78d6bf2dbde3be53634e232d52a793b7778affffffff162f29721e93b2c9de6629fffbe68596e94b26703923, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7e2f80300a4c81543e324e9c8973bbb6f16599c3d337ee82aed816624843f370, 264'h0080a807e920deaebaf3c3247010cb3c91cfce21b0d5ad695177d934ee5a7f7cbe},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{334, 1'b1, 512'h2b88c2f7b3ffbf92cf6698268ef14cba56c268701a73b30436de1465b85a572363de2fbe10e2beffffffff9b6ad94f832c537e1e40dfd29f836574fecb7dd074, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00de12eb33b717fd887fd684a64af9439a27ee83b28ac5751772249e600856b59e, 264'h008dca367bd7bc83709f25b0fc4e1f4a0e7e747be0b8a2977aabd25750a0ba60c2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{335, 1'b1, 512'h4e29d13bd24e9f13d5e31ac769469a23d44278a67b110f7bab6095667a3a5180bc8124849e31af47ffffffff94e438c9abcb1301833210026c068417d2da4b20, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00dee112ed7000c0776ba4fab09f439a844addb86c5046223397498ad72d059de4, 256'h7039b715851e4b386ea15e9bb0899ca21a4e6f4ecbbce4f706d29274806400b6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{336, 1'b1, 512'h5199a888f66bdde1285c6e1d75e11ca4a6fa67ceafbf32d81894eb60ba36c4786868dcb1384710d5d2ffffffff3d60d7798468aacd9f552c97fa4600343889c9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009d01032d95cac596e7df6c75965c3669f29cb8e58cc9a933bc5d60c1a97e946e, 256'h1cf2ce39df73cc734bb4180ef09de883bad7c8d82ab1a5861d265b48aa195bb6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{337, 1'b1, 512'h7692bad59be557b4e1db6cf148e5f0ff3c273d29d9017b90c8c26236cf78465b335a40716400ae0aaa34ffffffffd68ebefa85c403e0a25dbfeda3354bcc2a84, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6f1513d12e2112ec4f396ef4ea38324102ec3c7fb63ee49f485cb421a07dce57, 264'h00a78fbd65b2582a4031c34c7a8c28f03f16ef2ba18e2da41ef173ee5a85af1fe3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{338, 1'b1, 512'hadf9dc5a02f2bf38df234e566f0b5ae3c8b5a20cecc2f8565bb8f756ba59b295004e2ed1807a1e579596ffffffffffac7657366f92a09ca3685510feb2182e3e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c3fb59671cb8c6db48bd51a667060428f75124b5e990af1e997fd636335072d5, 264'h00c797e7245cfc8d98bca3ae1f4239b88684cadeda2c628f09ae61053eeb683771},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{339, 1'b1, 512'hf9db531c8bd06c7272a9ae2de6b4cac8e0281438eac5689c7f763241db7b88b4a6c71d53a3d03222f6195dffffffff0b690ef5a310f733b13a1bda4fe964a38e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e8b5b3f3443d59d7521d093884486e7a6732e275ec13313bd4d178f28128e075, 264'h00d299b062928e5f058c705acc3c62f24128ec703c28288b0d294216370cad69b0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{340, 1'b1, 512'h273f59b9ed631e0fc10467687508d817c2229d48e45efa2a6783290c6ab048c048a882eef2730e7456b3d4b6ffffffff0369568d9ede46d524123c6cdf78afb6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ce43218d44e113ec38d5cbcf402f3dbfa87d58826a760f0bf2c88f11981f7719, 256'h648f3ed0d1b76dec5437cb685dda7a1512ef07f4eb078dc50e418efeb1af8849},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{341, 1'b1, 512'he6ded1492cb08b685e2c14f2f11d4bb2fe1601c47019cdd5bb3a42aadbb88f1335fe76ecf455cde30b30e18d35ffffffff921892b8870a2d1248dcd97ed5449f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fdc99047865eeffcb69f8b8728a008e31f9f6ba78f698fae62b71cce79501888, 264'h00f06612f593873a13459695a5c4cb504acc2a8c56179b68553e60f2319c905b4e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{342, 1'b1, 512'hef9ce8e0e84c667ba940ccb1d3317daddea8b9888a2ef5b718605aeff060c7140522f73cdb7670b0e055a2646509ffffffff81c895857965435d4c4421eaaee8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h256e5c4f4cd121e2dee1987be7b241b6e91f90d483210aab9a4b367db5613174, 264'h00f75060db4bd6cd52bb8e6aa94f7ab68488a638873515787ec0d7e61bad58ab7f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{343, 1'b1, 512'h388b354799942c6595ba49bc6bf8e7ca5c06c6ae8015c0f58e69192d96cc60e30696c1284ba98c1b22c5c7f23bf8e0ffffffff15f579e355c7258262f0fdfdfb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c7a269986b6ad540dd30e620d1606e3267935c7fd5551b3311fd4e840510c248, 264'h008db7c8c464109cf0edb89357e663de6e882b6f5906adde6d58575ce0a2cce257},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{344, 1'b1, 512'hc6bf307fea8c2799ef482911ac86779072e5757f934a3671ad8c5a9e372bb2ec8d318ee3bd0cc4460f9050c937a3409cffffffff81c81c22e9468fd07ec09f55, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0bea324758ea80ed4a0a56f7d836fc73bf196e43fbc59d953f0ce34abba57b22, 264'h00f04027248e83bd48fb1571291ca1a5f088eb3e89f00904d71b9ea8d6677f7893},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{345, 1'b1, 512'hf5f21b002be6b7b3a605b3bcc5a3a12aa0b905565d958028fb8c44d8e5182b6ea4beafe63cbdd96daef63b98ae46ff91bfffffffff3ffcdb29cde67329851fd7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5b53c96d7a195f02cfac2d155aa7e132fbc35d59afb080f649dc13056248addf, 256'h2b157db2154bd5dc0ef2fc6eecd867fabdc633d2ca683a48f3f9095745351aa6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{346, 1'b1, 512'hd88d68932ee321d611334d87de84ef4240025f9d0c8f11bd9aaea2e7729ad87ab0ee66d229b2eb78221050b375a54bd698a2ffffffff0967dbcb983a8f09417c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h24174a81d221a4bfd8978f312acec4dacc4f08f8f8cdf29b2024bad2177758df, 256'h73fc1bf3388009e3219cf4c7e62e4aeaffc1b9614b2831405a01403c86936452},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{347, 1'b1, 512'h611df311628ef69305da2acf952b7289eaabbf389dae756f08c459819db39b7133f02dd126e0442f19bce8ee83cbaabdcd974cffffffffb7195ff14e2d445864, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5de7e80ce3137f5705d23397197c86e7749e5e682104f13beb5a6365a63780ea, 264'h00f3da2bfd6442638da60201be68fe2ad206365af9e40c4c1531cd3a05db1ad3c6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{348, 1'b1, 512'h4f34828f9520f17da9e588884a26df5ab85e8456184bb19001abc926a180c32a112ba4164e81d69b8fdaaf3c60619a7d1a5840b6ffffffff8748db5ab09c4a64, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00dcdc28f81ff5ed91fa15f15fc4f1d38f9cddfc3df65bb2d3a55582faf7c0910d, 256'h515b7759a130d667eff7ff3167c305cca101be3a07945fd7cb6a1359c16db678},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{349, 1'b1, 512'h4a3d25b54b17b001046f323462e30475caa0fe686e8fa4eaa3b0cbf604de9812e2cb4eafbbe44222356c1e1702c09078e7df08dc98ffffffffff06067e01ce41, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7407261c978018cc6e92a340de80edd3044a6e7116eb9fa9b022a2aeb318c65e, 264'h00bb5826953e0b85ad69745249f69507765a93f82198bca1e4475fd5de7dfb15ca},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{350, 1'b1, 512'h6a763ddd1f348cae57162f918abd67d536a03431ed29721e179403366c3fe64f1083d4a64cb7a9fddc7c5a3487675be4078be3b484ffffffff2d5a70dd12c49f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3962520ea2ef01cba7d5135117a7fcb5ab120b28baf6e31de2e6ec9993d8d5bc, 256'h2583659fbdf83399309bddc89ea5f39fe22187671f3149d94f96fa234a6013db},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{351, 1'b1, 512'h0844602883dbcf60972c8b943b5ea020ccb0d19c82eb86cb18d4225a79f97279539214d6e3df6ba6af165c9cd95b8b67a36b39bbd101ffffffff5a9aa9794dd2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00bec3ea35844452bb739d92b20882e5b672dc6eff323cd31d1a2db37db93791e8, 264'h008ef77b3c709d60b9d5d998f81d3f72c466fd7bb99c681ae8bc9c580db1f7c213},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{352, 1'b1, 512'h73672c1037e14e2ed10a0928e8938944667e83879d16f2688f2fe0087494b9f496471dd4e27f5cfddfc4b5efc4e7fcd511d2f67ea879f2ffffffffaebc4501e4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b8fbdfedee5376cfc9177d96c45e003f90b7367aa40cf37d63e483bfaa4be951, 256'h4dcacdfbe41df7899382607489bb75422f3eb67822890ea3bbfd80cd456fc127},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{353, 1'b1, 512'h1c28cbb7dcfe2b79763ccf8ebcb7939ea373f7751d8b3965fdcd8b62e8360f619321855d0fe872fcbb3509f48c195d96b1d765983c695686ffffffff51d7cbd7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00df228c1a8bb3684b7ffa2e3f777643c369e1bc2299d66a66c8ed27a4ed59b783, 256'h47314aaf3629a0de02313df06c0cb363e4e019aafd20ec06be63b7b4c21538ed},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{354, 1'b1, 512'h823e30e3f8bce86e5790d073d931eed5a7ab1f52fdaa4a2522831c73dff05fdcc91829a51c8c0c97c24def713b52643ab17a700ddfa0988740ffffffffca2992, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h528746b280d8a0e54851cb99894afc01ce24cff7edd60116e3d8dae42adb4961, 256'h4eb264629e5cf4aba77e05c54774bd0cf20b057142a1ac2103099d664c2c5dee},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{355, 1'b1, 512'hf2104bf641a8b485448e73c4b7de7fc4ec1d3e06eae0f264dbdadb0d514a7aa2ff1567a80e8156c2bd97579eb1467c0efacf0fdd1166e87838a2ffffffffc8e9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h44c391f82cf5eeb80f87c347a5bfe461c49fd8779311e237abc05b19f6aed093, 264'h00866853619339b716092df4466aa0cc9e6256fb7e18a79854b60ccc534bb6df10},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{356, 1'b1, 512'h3db47a2cad8a1c43f31ee677cef231cda0f3853901676c1732771602ccdcc294a38fb8df77d5e6e5737d4c8e05953aeb81edb39a25931717b3c154ffffffff9d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h03d127a6f72465bd1c02109f9605202b246763097c756235d8f8a26848eb609c, 264'h0083d551427f31b9572b61180cf18bc85c20306c0de2c39d00430b3fc91dc50c6b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{357, 1'b1, 512'h6becb022ae22ffc4efd852cec1259abcbd9936403db48920bab66dff9bd34bd1ba5c30d1e8752af80d13d9304dfb864e834181cff7e8be9467cc3617ffffffff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5044ef2362c8e6c32fc14584b0751eda8e8e8901d9382354040d2615d9cc07c1, 264'h00dd16765911dce7a7ae5f3b64b3ce3a5e12e548784597dc0a379f7bb8f4fca879},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{358, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ce645f0f1ccb63844e54bd7603a4280ea065e3c147d26e73cfbe58c6116b0cf1, 256'h40ccc23188aa20453d7f95d33868f247b3d77c516b70e4c351b48ca2ebef0027},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{359, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0fa36769835d1d215f156d5e82bed2fa76aab134bdb1d3bd40975faf5ac19cc6, 264'h00e67d675a8f0dc4760b3f8fbe0f0853a80b58af8dd2c4a41afbf9cb0c72d016ca, 136'h014551231950b75fc4402da1722fc9baeb, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=136b(17B), s=264b(33B)
  '{360, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0fa36769835d1d215f156d5e82bed2fa76aab134bdb1d3bd40975faf5ac19cc6, 264'h00e67d675a8f0dc4760b3f8fbe0f0853a80b58af8dd2c4a41afbf9cb0c72d016ca, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2c, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{361, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2f1db0895a8d615779a38ddcbeacad9458f35688b587abeeda1cb5a891e954a5, 264'h00b591478e3b81f5881dd71f93b811130a67ea697f452faccd5c5117fac15f5f93, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{362, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h462155174b64dd050601b6d7c2297251815d413e26c9b91d123536e76fd3fb13, 256'h5f0a20f86528dff246ecc71d5d005b2935e4d8e0b076fd6792d4a2b3fd2b7bb9, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3e9a7582886089c62fb840cf3b83061cd1cff3ae4341808bb5bdee6191174177},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{363, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h008e89e0fff2d768c7c139b22b90aa66b24b3b1ced4345c469e439b2c80d6fed08, 256'h4eb9ca1486ff3411db46590f78008d6d6a0a9cf9cf36b2bef833407af5bc883e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h24238e70b431b1a64efdf9032669939d4b77f249503fc6905feb7540dea3e6d2},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{364, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00f4c2d7df7ca616bce49212e47ed112106445f47cf114782626740d37e1c596df, 256'h1088b19bcaf0d10609a46bbdfd626a83d13e62d405775ae3941755b278a443c0, 8'h01, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{365, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h43053fa57436a0b26f0f887b2403ccd9d18f14b7866e1da593835e93cd103a15, 256'h6039d7ccf6c355ac94ed59225aab8a5aa190c89c422f80e71246b998818ecd54, 8'h01, 8'h02},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{366, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h009b27e4409c49abe9d8d1b90edc64367daedb43d68a41c501032dba5d73ef1021, 256'h0cd42cc8488eb0588680b94e934ff744f4e6cb079737beb5eeabbe56fd11a7bb, 8'h01, 8'h03},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{367, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h009b27e4409c49abe9d8d1b90edc64367daedb43d68a41c501032dba5d73ef1021, 256'h0cd42cc8488eb0588680b94e934ff744f4e6cb079737beb5eeabbe56fd11a7bb, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h03},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=8b(1B)
  '{368, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6e3f0e1b05e5bed7e8a1c8de7b8a1273673731151e3a04ddc83e18c98d842943, 264'h00cf1d41058a6b7272a014c6caff94db3f0233e0f21cc101ea159ab14bc8483745, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd04917c8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{369, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h06b2c1b72f12846bbcceda68183372d3f05ec591c43569361646f5916a00a720, 256'h2282d15b70f19db914c6fdd8faf15ab90ced3bd4c3f59a247be41610497594c6, 16'h0101, 264'h00c58b162c58b162c58b162c58b162c58a1b242973853e16db75c8a1a71da4d39d},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=16b(2B), s=264b(33B)
  '{370, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h4e61226e0b1c1e5a40767956c7b530eace83d550038e32bd14c5258c48c939fd, 256'h57d069215ea210b386820a2d426fc711862bcfb34c7deaaed404d17692892cc4, 56'h2d9b4d347952cc, 264'h00fcbc5103d0da267477d1791461cf2aa44bf9d43198f79507bd8779d69a13108e},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=56b(7B), s=264b(33B)
  '{371, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00cf259a52f769eecab5071c0b4676bc4cc474474b74675fe8bd1660df5b70ce1b, 256'h722f774a601a61f2e8e364477b0ccea457b76977ab300139c4ee0e1fbb7fe8f9, 104'h1033e67e37b32b445580bf4efc, 264'h00906f906f906f906f906f906f906f906ed8e426f7b1968c35a204236a579723d2},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=104b(13B), s=264b(33B)
  '{372, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h67ba78328cffa6eb3f7119096adf17e3fca6b2da966c03bc66174c2984a1d553, 264'h009abdde7989d6f5083187261393a6e162eb508ae62749e41caf55b2be14d9a960, 16'h0101, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=16b(2B), s=256b(32B)
  '{373, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h008f8c5fdf711aff7ddc807c4308a132b1099e3e95dabf803ca29283dd41b09055, 264'h008f60c71b4a813e7b4364b0a7260765042d3696a9580548f585be12633ac3b824, 104'h062522bbd3ecbe7c39e93e7c26, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=104b(13B), s=256b(32B)
  '{374, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00fb78c45f16de9b4e098ddc9ef6eb340b055a6a49c438b87bf7969dc24f7967dd, 256'h2af9ebaba55b6713e06e9df9e42b79ea9364405ebab1199ea230ae38ec83b91a, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd03640c1, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{375, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b7b91538786272e70a603cfc80c52f87f057a369149848dbc865a8d2f445ec26, 264'h00bd90ba8844f58db6744b5f31a470e59ebfee1891be36ee65b18ba172e5eaf943, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{376, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b7b91538786272e70a603cfc80c52f87f057a369149848dbc865a8d2f445ec26, 264'h00bd90ba8844f58db6744b5f31a470e59ebfee1891be36ee65b18ba172e5eaf943, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{377, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h009c0c462658f6493295775ed99348db5895ae8471c819a1ed9ae1b5180397f08f, 264'h00f386d14d6e56758d1dafa50755af4fe079233c139436abf61a9208f8b7f893af, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{378, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h0089e63127c97dd4cb19fb802f22229decd0d852639b3d982b2589817a7e520049, 264'h00e1fd70b15e5e5d3ea4ab748903ca891ab3964ff4d7bf48b17c6007957a5e2021, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{379, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00eb89c838542537c3f530b6e8bc62d1e6284ed4e9b8c6aea96e82970d8abdefff, 256'h58cae0df61874d30c2afa05c8a703800ac80564397688b19a5149f65054b138f, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a1},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{380, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h72bdb42d379cd807e8dcdd597e5c68c464ecb4211ee885f7210e55ff52e93688, 256'h34231f3921839c8a3a2cc7ff5964f1f79c77f2c8813e2659684ee1d8bf7125c0, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{381, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h57cf2c69876d8a9822a6b796492aa889c39fa1371fc730c5a15532ac4aa197b3, 264'h008c936d0041821e1ca81df3f1fd0a495c0c8974a81fb41cec4622cc1bfcccf3d2, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 264'h00cbd2518ae59c5c357e7630cbd4c4cb1410897703e7663f19fe1289497bee4f7e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{382, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0a7413800a6571b03100d9f327c68a89aaaef2e7ff922b0a0aa95e39a082c4fb, 256'h37466eb04ed38187bedfd767de7c45416577bca4bd961de3d8890bea3409f697, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{383, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h7e27893adb379d40a61668ad660edc256004bbfc12d55889fbd5121eac56a06e, 264'h009a36f42598db7d643842a72562fe6d86ddc38623830e42a17d444d44a2472b5f, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 264'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa9d1c9e899ca306ad27fe1945de0242b89},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{384, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h3b65f40a248d91a7e6377bfb5989f47d562bdaaf364ea982830f61b71957bda5, 264'h00e42108c5d388f2e173210f867633167eb0f5cbc693aa7bb9223ae8f1aaa26983, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00bc0f3a2708cbe1438083451163be66f80a810a900cd135ddc076db7451917c17},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{385, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0585249ff4a3acbb996eed6f17a70a7b83a6dfe96e80edc0cd4cc7594e806d59, 264'h00b7576508dbb4eab123e0ed688a9e6625d056c7ad8134776252728dcae375cd84, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h62bf43ba34e73cc3c8922f26d64e3bf882f12dcc06e0b30c8363efa6badcff55},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{386, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00dd6ba66855e37b7fc91ad160bc4a7c5089f8633ac0e12298a6aba34db680e16b, 256'h798f5573bd93756e39dd635d9c5f8e876364445a1c9a43f2918beb9137ba3b92, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h39422623a4386033ccfa96ad4f8228fb88ac9364ae8b3cd0715ee188c467572c},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{387, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00ce2d8a8432670515b2133689d96e7369decfe994c87e39a28e5636897a360f2a, 264'h00ba43f7fa77feba76de9634b6adfde47fb16f70b790bc9a1a5065ef16f6fd2467, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6233bcf8558bae02cbd2518ae59c5c3501ab620efcbd7b40d8dd1f7288ff5dac},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{388, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6cefd89c949069c4ef5fefd20512a6fde92e08a2dfc408694a05d2a974bd0284, 264'h00ae4769496c219a59383a7fd6dc1e0690c25506264b0088e0362897e0da59103a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3bcf8558bae02cbd2518ae59c5c357e7170b54262d04bee3a9fcee6e38e84e1d},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{389, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h33a6ee1a121ccab25b00fbecc860be15641a5baa4b4beb35d9a6dad35a1691fa, 256'h36ba2323e463d684219a1bd15c5eb304878d82d1da113c52c7663cfae3f5751a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h779f0ab175c0597a4a315cb38b86afce2e16a84c5a097dc753f9dcdc71d09c3a},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{390, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00a2d2e9810bf8f988af6cdf111f2f15062900d2ce06bb72c9c1dd1ca90d69c58c, 256'h36c24fbc1323359ffc3d7cfdd66451dd3e950ad97cc7f1ddedf30e3aa4425c0f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h558bae02cbd2518ae59c5c357e7630cb680f5a3ee98045977a021c9091920d08},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{391, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00e93d658ec3a9418daed0ee219d18180d0684fd676ed24f693bcdeb7e358ec44d, 256'h6914850bd227eeb22bf22a02c3bfd628c769b0f0e50040b50fd3aaa324a1d4ce, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h19ffa32fd51fb796c6154167347b7773d9058ddb148fdaef8c287fef848f2f7b},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{392, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00ebe7e1278636290cb09c7d4554c71c117337d2ed40c77789433c27eaf4d4bc32, 256'h73025752ca492238b622884c9fe287ce3723ae04ebfaa53505e14b8e86c5dbac, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3d180992c1a38ddfd49ecf3d1813b0b195c69b06bbd41cf101fe40dac9c9e6ba},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{393, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00d1150530bac21e35524ff9e1b7d00731401072d591e696a17bb388b4d7e5ca19, 264'h00bcc66bce3fc176d2da4a2cb954c836bf9b81f1913230ba99ea6e5054073ddf6f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00d39813c8e58536460cbfac4b0fa028e60d5d45c13612d79f9964a58cb33be185},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{394, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h5233a1deddbbdc29c0994fd43ceda3b020b35c465e02d1c12fd29017306be87b, 264'h00c31db5c0e32fbd3f045664acf088014a1116eb3379f24886b3a13f009628df42, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00e9fcbcae7e1d744cf6bf4ca0d8573312a131fcb3b90eb26bed6c7f6ba908ab53},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{395, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00a160ab41fd3fe7d088ee874c8b82d8ae97c8ed99467579d01b97bade23ec46a6, 264'h00ae709a088bcbc72342996efeed0e913f8a5dd8c8878b1caec5c9e057e35d5cfe, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h21f862ec7b9a0f5e3fbe5d774e20cc835816e92b513bb52effadc18c3f526295},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{396, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1d915ecbbf4c25bbc0d2216db6d1a3da8f80058653a24885494aff88fe1599fc, 264'h008816898d958fa5431bb557d17b6b1b520c3fbdab6bc5984109d1468b6cc141f0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h43f0c5d8f7341ebc7f7cbaee9c419906b02dd256a2776a5dff5b83187ea4c52a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{397, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h009598101f8704e2dd0e889ecab9ffe7a5e7536f3ee60d5f05111ce6f5a4ca0405, 264'h00c4c39bbca34c6a687c46a6ddff65e81d0a9a78a8c104f91ea6636a7c8ea6819a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h65e928c572ce2e1abf3b1865ea62658a0844bb81f3b31f8cff0944a4bdf727bf},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{398, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h59ee9e0a000baefbe3fb59ea61d7370df77c58dee9d829b6c5e89faae019951b, 264'h00bf61a756c7a30d049bd37010b7b1c25670d4ddb6ceb8f1d7c7d449e393465959, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h1ca11311d21c3019e67d4b56a7c1147dc45649b257459e6838af70c46233ab96},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{399, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00d1f1ddd12c710d7c35617a0ed2fc35f4d09888f17034a47fe0a78415858e66a2, 256'h5fcda6abedc3a58ffc55bc5d9f320c60eb6b4c9a22833e13511b2e140ef14057, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00d55555555555555555555555555555547c74934474db157d2a8c3f088aced62a},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{400, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h3c9a5007f19ec624a73ce75fb61ab3e16736d519ee36381497f24bfd3bb691b5, 256'h34b42b0134e17222eff05f3b5477323a3224310b108c4a8fc9b17833128cb822, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00c1777c8853938e536213c02464a936000ba1e21c0fc62075d46c624e23b52f31},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{401, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00f7a2f1027241c8514b2be7097a3eb5b208e8ffd09a700e5d72fc3af6964b3bbf, 256'h08318a9043d959a8fc8bafa5d403d3490e4e45d9b1e156ff3e2aee38ece66e88, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h30bbb794db588363b40679f6c182a50d3ce9679acdd3ffbe36d7813dacbdc818},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{402, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00e58d8aba787d54ffcbe530c5ba5955f54e286d31f1a7558dce8924000d7a1b96, 264'h00f5acbdf479b313380325edbbadbc6287e08e98cc86e2ba8339873724437ce813, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2c37fd995622c4fb7fffffffffffffffc7cee745110cb45ab558ed7c90c15a2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{403, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h167df009cec2efd44991a523dc2fd4a13e4de3e76390382d4c1088593f33da65, 264'h00838f62138f2ed73fbc7be316ba5b6a79a4768fd1f4ea07df9eb0eeeef988ab73, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h7fd995622c4fb7ffffffffffffffffff5d883ffab5b32652ccdcaa290fccb97d},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{404, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h01a3a8df8aee278aa306844d60d9c5113e596d66cc92a3566ab0797cd0163825, 248'h62494573ddc9a21706030fd795708b3fe0d0f224ac01e5957ad0d11d6ee265, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00ffb32ac4589f6ffffffffffffffffffebb107ff56b664ca599b954521f9972fa},  // lens: hash=512b(64B), x=256b(32B), y=248b(31B), r=256b(32B), s=264b(33B)
  '{405, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00d6d0f45dbfa12ab4ea5b29a848c71923d1ecb57b148ec1c969b43662a18d00f9, 264'h0088c2728d21508a421af6b612a4433c4b7c97f55dc12b24db2cf6cb7fada43f15, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5622c4fb7fffffffffffffffffffffff928a8f1c7ac7bec1808b9f61c01ec327},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{406, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h69214198388da2a0d1a0c9464c6eb3731ad44e27287c17cd24bf73c3ada67c2a, 256'h48dfabbfa5d9127fec9fb7986fb386cb5c7ebe3f609d95e71a70ad7f83334584, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h44104104104104104104104104104103b87853fd3b7d3f8e175125b4382f25ed},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{407, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h0084672e2de042df2668775733c9b0cc716edd7d7534eb859279316ec5186d7733, 264'h00badc81e933abf3d4ce75fae00d1a47b30d69de8754666a294b4c925807dc3ecc, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2739ce739ce739ce739ce739ce739ce705560298d1f2f08dc419ac273a5b54d9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{408, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00c9be9c1906a73789a9af1a677f60dd4163c5fa06c7f45c0993a63051aa0c0f30, 256'h3205debee5dc413e4abb3e1f6af550ac64c41b97e425cc2efa2a833c2ee72221, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00b777777777777777777777777777777688e6a1fe808a97a348671222ff16b863},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{409, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h026794f7b5a84849f41141c68d3248f9c90c4de7edad4fb8f446e3076ffb7962, 264'h00c98e7b67192296efe04379c6a40280b4f113876981b44b73bb676a881f398790, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6492492492492492492492492492492406dd3a19b8d5fb875235963c593bd2d3},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{410, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h18bd65dd46f8c0e326553be55e5e234bb43188ac1fddb37003d12f091aa7a1b9, 264'h00e9c00a03e4d5452ba9a607951d4e4d8a7391a952109d96599266d1e2d9ab2199, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00955555555555555555555555555555547c74934474db157d2a8c3f088aced62c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{411, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b86ae764f2f95eb9331af538fa516fd78435794ebb244c090c6d6b286750f94c, 264'h00f3712f767495a10f2e81350662af3ba09defa2e0e6f27eceea35513032dafb61, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa3e3a49a23a6d8abe95461f8445676b17},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{412, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00e045cc5a9414e45e63f1b08648e20e229a9950ab56ec304e1b907989e81af2bf, 256'h21e52db489853dc470713aaecd6aadc7bfd8504a9c82d0243f6e774600b5ea0a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00bffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364143},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{413, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h37e377faea8a867f494bb402032c70c12af6fd57feb3866bfc5a5fc1d0a909f0, 256'h08dcbc53fd41b67073a4e71a81f3fe578da4d5add0d698041a9b7f38a9a19bff, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h185ddbca6dac41b1da033cfb60c152869e74b3cd66e9ffdf1b6bc09ed65ee40c},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{414, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h09a33110676e4a4f8a977150a7be291e0a269cae9678710b1d87f8068b0fe961, 256'h043a6f64e86278a656a39e4468b3472597afb2dcd930ccba1b1ea2c988c13450, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 264'h00c55205f423611c7e96615bcc20141945fde24bbce956d49cd43e14ab4cef3659},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{415, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h09a33110676e4a4f8a977150a7be291e0a269cae9678710b1d87f8068b0fe961, 264'h00fbc5909b179d8759a95c61bb974cb8da68504d2326cf3345e4e15d35773ec7df, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 264'h00c55205f423611c7e96615bcc20141945fde24bbce956d49cd43e14ab4cef3659},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{416, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b7021faebf4081a63094d8ea78ca2004d02a303bbf363470ea4a649b08c1995b, 264'h00de5efba25c9d2f490f181e16795d5c75f83b5c11c81d67ede2ea8df81d970cef, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0, 256'h33333333333333333333333333333332f222f8faefdb533f265d461c29a47373},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{417, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h4de024ff2abe7af94fb5e9f53c87d4b4bf1c5447c7c39a9280839f12e52e38d8, 256'h3ce6941fc329978e794abf91a25e83463f8eabcf106d76d4dcd92c0ae05493f3, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{418, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h425e137c5fe08e842c3bcc4efbb6c4bca89edda8d6beb130e14899de2f20b74b, 264'h00b1af66ef5baead32e7892160deddcb57f43503104dbc331fa20a8de376e5bd17, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 264'h00b6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{419, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6c63d82f22bbeb1bd1c8eba4c680ae17dc2b4d196a0da0e191dc79fefd85e367, 264'h00a883018fb8d160ca01d17234fa0b060a619215ccb9dfea629d6bf92cfd8ed34b, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 264'h0099999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{420, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00dbf77c566f7483d7407f0095b8b468efdf85b7476e614b8658bcf5e71e6fd588, 256'h413b50407df0def01b8fcba5621028a6cb0972831c893e3d3c20065b75a8e8e6, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{421, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00a7967bfb54cfbd8d13492b9ac421d967d7c4b0a3b18efb6408a424914789c8ef, 264'h0090969628e6553898c978ba48eb852714f9e220e5e93cada91478ce1af8948fd8, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{422, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h325fd7ab7bc8cd7d859687937a90083f1b46776c2b8fdf4ce2bd9e2e808c68b1, 264'h00bb0d689ca6f542c094c99c71918f5455c7608514149148470494e05aa4ff6110, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{423, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00d637dc3c63060a0b21b80d6dc8a97ab6a543c21c18cb5e5c63ad80c3b86050fb, 256'h1d68bb9b9c36ade49ddd84c7fa3ae5c70f45549592ee03a23a490a891cc70ebb, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{424, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6bc87ce6047a3164be15ad781ef32d12bad8caaef7707ac3e15a53ed75efc90c, 264'h008eee286e2ac0c8f9f6f0350b8bba94b6c5bfade87ba211adc0cad5f3818091e0, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{425, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00dac247040488bec28dc3ec9a81a990701f45c0ba4bb6e22573da400efaa65e2e, 256'h7de375486e1757b6c7b4269bee423edb84c7f4b333c1557b5ddfba0dd983ccf3, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h0099999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{426, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1d4d073190b327ab4e4f5ace8d8c8b68e100fd2565a1a4c4610bca309fe6a9c3, 264'h00e274a19b41e496b0832e9e42f5229fc000706c966d2557f3441d323d8faca129, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{427, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h274ba8da21e4ed44e218320daa103f0d4227bb351b67d84ad2628629b82fa827, 256'h4c90d1dcfe55fe7ee66571ff4526c755cac8c8ed16b01c4db830b7dd9deae749, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{428, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b45406f951d31975e953ac11c25c238046a7975dd2fbb38d890913c1c8b451cb, 264'h00cae0be688e6e400a9265bd9a59ba1047e164306ef6cd358bc0ff00e9e027e957, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{429, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{430, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 264'h00cbd2518ae59c5c357e7630cbd4c4cb1410897703e7663f19fe1289497bee4f7e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{431, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{432, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 264'h00cbd2518ae59c5c357e7630cbd4c4cb1410897703e7663f19fe1289497bee4f7e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{433, 1'b1, 512'ha69f73cca23a9ac5c8b567dc185a756e97c982164fe25859e0d1dcc1475c80a615b2123af1f5f94c11e3e9402c3ac558f500199d95b6d3e301758586281dcd26, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h22bb0000e9648a0ee659f9b6a9ab6513dc90ab968ec49d3953f64c82bddc8520, 256'h4aa0dfd047b0786e118231eff7e86311487ec9d1bc84aaef1f736f4178c288f9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{434, 1'b1, 512'h86fe1b4ea7ac8e339d04e40087534c61e245dd4a0c22754a0622642bba56de900b2d431e859a36b1a5ff71aee560522eb0d3251e018c2cb6a10b82031cfd37f2, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 264'h00855b60549e0d84ed3959ab2800eee0cbc9a2cecae2e510ed51e9f27975cdcc4e, 264'h00c60dcc80a3dcce9911cb9cfba123b6a6f85d20ab695a9ee7d46e0bd9eeb337f9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{435, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h5cd73aa58188658ea513f8ecf0d9e2da9eb5d6bcc7cbadcd6a4a8e0cba5176de, 264'h00a9f090bb5d3fcf5b7fa7e16d287718773f5f4ba0973b329a3788cd45b4bd3765},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{436, 1'b1, 512'h7d795fe6a97761d89b35f64e09555951f6ec2a669a9fa03481c100ae158f183e2171e142437d2c3a42352108a22a7e3d797beaf6c3075db419b6f4acca479c83, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h7f9eebad2a323f8346445d1e2fcde47aba4c96ad4686172bebcffaa604e8dbe3, 264'h00ec09d731e58e3a337ea03ab72612b1f801b88eac571bd3a031250ac6f2e34fda},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{437, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 264'h00c28ad156fe809ed36dc80812ae2f32d84dbbfbb9400123305c332551c4f10d39, 264'h00fc5b95b0c7fbc2e7cc4ec1bf01020f8050260ce2ca45c3bf5b64a7b2aeeface9},  // lens: hash=512b(64B), x=256b(32B), y=232b(29B), r=264b(33B), s=264b(33B)
  '{438, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 264'h00a36bfde0f5e23f6e3b3d6cc80ede3d9e4ea1c2cb9337221388f70aa52dec5e53, 264'h00c27e1db10d29720a120c2625c7e0756790200b2d9bcceb170a1356e1d5477e3c},  // lens: hash=512b(64B), x=256b(32B), y=232b(29B), r=264b(33B), s=264b(33B)
  '{439, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 264'h00818dee9730f01b3f525daa9cc0d5423b0c4af0414c647b6e0bc88546db9c0d75, 256'h61c16a90de1dbb1ab1e3c7917e891632f557f493b4106f225517ef186abc0ff9},  // lens: hash=512b(64B), x=256b(32B), y=232b(29B), r=264b(33B), s=256b(32B)
  '{440, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h53cc0edfc688e3d264ed4755f9cf006418e16e24dc978453a6ef14fbecff617f, 256'h24694c00d38c13259973aa6db88adf7cc49b5673e628b3c65e7fe06f2665db86},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{441, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 264'h00cacd14406211ed85d8de1b50e167f59dec688574524c6fc1762c9268214e3bba, 256'h289cf8949f717626c25833a0a159d63d77d022b48e161007464f59f5072df8a7},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{442, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 264'h00c1a4c9d1feef48045813d911f6abb188502e06d26b34194f2deaa356e578a769, 256'h4063d3367b2bab52bf9fbc4cd3f670667569ccb1cfb05a7c7c156622ba593d45},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{443, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h5af5683467b4cb3d68bd168c5fe229a07b7eb1de2f92b8a9743fb46c3691872a, 256'h4cbe35cbe66805729e907462169c13b5c4feb497aab658774bec1ecd7bd8863c},  // lens: hash=512b(64B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{444, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h051e5f825a5c29f92a108a3ddcdcbf7ffce37ab32915985978512e89a2a83b0c, 256'h6340ac187077a7fb4373537b4595a39299ad0ba351db23bcae9176125c61eded},  // lens: hash=512b(64B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{445, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h34e28decbf74abd30f55155ee2ff96f621066001a853acef916cdb39a7d07b40, 264'h0087561a96167016fb7dd6f3c7259f8c563f2144332ebb9a48e93b9512d3bf5392},  // lens: hash=512b(64B), x=232b(29B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{446, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 264'h00cafded1bc98a4bdfe76e1df9ab75342a7fed16b0c1688a2e744d871b9404be14, 264'h00a11fcb57d1212068afed86a37e7291aa02061e75b883e9b9a7af3a52e81f5033},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{447, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'h254f9541aebd4fca9ce7136fa8e6ed6367778afedf36201779b0ea6a61a82f3b, 256'h38668103eebca5e786e05dfffd8b9f1d87d4a1558b1cdfc0eeb98a606ab654c6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{448, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 264'h00f998e8322b2a1101bbdf9b8b80bc147e5225632cdb6b1a8c4c4c25c29cd3319d, 264'h00ee6b3e7b59621fd62b3253ef646ad7cd4a4d53dd11372038b0b314ced0e2e5a9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{449, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'h0c426a3f25f5d0250928ac4e5ea03cf949d34444283ac18a49ec638a2a6ea4c5, 256'h09f0df2fe78f8ce301057c734cf3c2505d7219775fb778758461360b168e2c8e},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{450, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'h1309ba742999ad66aef104cc140246bc576bd14acc6bb0be728577e49f4f8ed5, 256'h31e29fedcab5999d66b27a4f4ffc950dcc8066fb7cdbad9a6362270c066a500a},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{451, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 264'h00cb565ebfd48044d17d2e241b7cd5fec6089e3d0bee83516b710f68d583ccd1c6, 256'h26d6d5a1f12ae063528e7e4b1a6a9c5c760af38f2828db9407c439484f2ae9c1},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{452, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 264'h00a6c419f478007ce4eb07cd8deb248b8d9d11e16c02364e18391ab934c6f3e91d, 256'h363ab461b8d40c864998a6dfa9c9c77419930b9336f0cd471b74786b09aba27b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{453, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 264'h00e22ab46f883c6ea58de97f982ffd3ef581749fe5568f8121761566509145b0c8, 264'h00fc4a53daf4122aa10b98a4d18c2e4920b37744447f0d843ff9ed1d79d482d73c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{454, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 264'h00921a16ea241e69c9d4f3bde6ba2cc7e10a27c9dfd8b92076d0a4a6d9f8ae0ab3, 256'h39b66ee2afd7db1099fee2cd8c69c9f1ea29047efacc1c6e8ee92e5a2244a40b}  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
};
`endif // WYCHERPROOF_SECP256K1_SHA3512_SV
