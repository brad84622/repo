`ifndef WYCHERPROOF_SECP224R1_SHA3224_SV
`define WYCHERPROOF_SECP224R1_SHA3224_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp224r1_sha3224;

localparam int TEST_VECTORS_SECP224R1_SHA3224_NUM = 252;

ecdsa_vector_secp224r1_sha3224 test_vectors_secp224r1_sha3224 [] = '{
  '{1, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 224'h56c80970d9a308a9f639ed199ac088f93ba9afd04c53f48e4fa88d3a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{2, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'hbdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{3, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 224'ha937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{4, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{94, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 248'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac158453760000, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=248b(31B), s=232b(29B)
  '{95, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 248'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d030000},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=248b(31B)
  '{99, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 248'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac158453760500, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=248b(31B), s=232b(29B)
  '{100, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 248'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d030500},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=248b(31B)
  '{115, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 0, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=0b(0B), s=232b(29B)
  '{116, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 0},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=0b(0B)
  '{119, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h02bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{120, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h02a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{121, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac158453f6, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{122, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d83},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{123, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac158453, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{124, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 224'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{125, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'hff00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=240b(30B), s=232b(29B)
  '{126, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 240'hff00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=240b(30B)
  '{129, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{130, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{131, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h01bdeb8edbcb30885c65bcb58d6ea1eba154c61a02d5e2fff171e07db3, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{132, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'hbdeb8edbcb30885c65bcb58d6ea3be5b93543986ae28ad66b9282939, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{133, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff4214712434cf77a39a434a72915d2b018bf2d63b3dfa2953ea7bac8a, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{134, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4214712434cf77a39a434a72915c41a46cabc67951d7529946d7d6c7, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{135, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hfe4214712434cf77a39a434a72915e145eab39e5fd2a1d000e8e1f824d, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{136, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h01bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{137, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4214712434cf77a39a434a72915d2b018bf2d63b3dfa2953ea7bac8a, 232'h00a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{138, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h01a937f68f265cf75609c612e6653da44c85c830abdb665dfc690fc740},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{139, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 224'ha937f68f265cf75609c612e6653f7706c456502fb3ac0b71b05772c6},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{140, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'hff56c80970d9a308a9f639ed199ac172565af0bf923876cb48f34c62fd},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{141, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'hfe56c80970d9a308a9f639ed199ac25bb37a37cf542499a20396f038c0},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{142, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 232'h01a937f68f265cf75609c612e6653e8da9a50f406dc78934b70cb39d03},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{143, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bdeb8edbcb30885c65bcb58d6ea2d4fe740d29c4c205d6ac15845376, 224'h56c80970d9a308a9f639ed199ac172565af0bf923876cb48f34c62fd},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{144, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{148, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{149, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{150, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{151, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{154, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{158, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{159, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{160, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{161, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{164, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{168, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{169, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{170, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{171, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{174, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{175, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{176, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{177, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{178, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{179, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{180, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{181, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{184, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{185, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{186, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{187, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{188, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{189, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{190, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{191, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{194, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{195, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{196, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{197, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{198, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{199, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{200, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{201, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{204, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{205, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{206, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{207, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{208, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{209, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{210, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{211, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{214, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{215, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{216, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'hff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{217, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{218, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{219, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{220, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{221, 1'b0, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{230, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 232'h00bd6b1d7ab97ac1b607c22e042ffcc0062c744160c958ad0b1943a944},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{231, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h476bab7a32e1f66958492deb681033dc135276f62d9265c7c7fddff4, 232'h00bcce78ad8017bb499490eb1bf00dd9f35b23b5e8bd03fe5bb09e3f5f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{232, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008355270aae4ef8dda33cdb3fad664dfb0124f6dcc0e79a9a7b6bb19f, 232'h00ec8d3e43977e2692ec27c702a6f349d4536d00cc017b55f325227da7},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{233, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6222915ddf6e69eaefce3ebda56ac501428b3d69b7b94c0e9ccf0010, 224'h5acbd1d130b50c08778175172a9d0d0e0e36b6a68c80af9aeae41b6f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{234, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b8e3edaf6aa9e6322e916ba1cd2bce6ce694ca8e8f9f999efe9cc07, 224'h793b8d557b98e504bf05b2a57b1fd1eaffb38eda30db7c5e8a559c93},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{235, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a8b78286f4b4ade20d7a8f7c1ce3c29d6616432eb99b34cf8a46d421, 224'h66b05e86c8a7e41fecb51047a7b8d7c4a6baf806e9d360f0c6715c6a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{236, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h33529fcafcd107596f846563605f0d9c479f5ac9498e325e034fd001, 224'h75e231e760bc10eb97901c2b8ccf908099ce7fc54472fcb419784d36},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{237, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d4514aa4da10577bf2974ff7f6e410e82f9267877b73631e0b336ecb, 232'h00936e3ddc7846ceebb4f9e8c262d014f8ec5ae90cebed2359b49aa559},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{238, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h65d35e97f9455bbc13c8ec28f8b8d13ab7327fe77c38b40f5b855c37, 232'h00a21cad033d04659bd2539e7838e8377b5b11f14d0c016616775586f1},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{239, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d444ef96649d01d2a47a9dd6210b45fffec0ed1a4cb7438e8cccf048, 232'h00a828341bea5c28b55097e77332dd7e303df789a2a67946de23dd3473},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{240, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h09463baa1c7630494a9ed5d64fa2fac19ac452b3142f8bf19f585574, 224'h3897d58b8aff942a074a583604b174ddeaf230d7cead58e74835d89d},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{241, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4c2ba44adbb44f6b0f57de21830870d5acfc68e03c8f35e1dda14cec, 224'h6aff00cd6417ac43c1ea7e107fcfada404b88f4a79a0d12df96ab028},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{242, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00dbbc41eea7c5c204388b7941cd19acc7a2eb38b8e848845bcdb4244d, 224'h7c4e411b930f26ffaa494d2522381ac86f38b37591d697d1229253cd},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{243, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h595b6900f6eb4494366219c35b40397ffdb3141bffb2d8d216f97973, 232'h00f53261795ddfb36ed4a83f783710f15a8f606cf9fb3f9ca1981f2605},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{244, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6a785a5bc1b857f7c10120d85f36d9d444a5bb6ed0991eac4a5a26a8, 232'h00eefa7d6774ee5851dd7f1c45d204fff4387ee126acbd56452d342439},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{245, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4e0f67b081cd6b87e3f4d792f1ccdd66e780d8028eaeb5c40047b615, 224'h14c42ea50c712c3fb7a0e18fe06b23822e9063f15bf2759dfc70383e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{246, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b16e31a9a07bed7d2adab9bfbf9fb8a279f6387791d229e79ff435c7, 224'h0cac45c70351a77cf2d0377601be4f7bbf5acddf0310f9e10b1c7022},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{247, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008753a04e4ce34ab8997df5f36934cd16368cb0f3e849890d74242acc, 232'h00d035d2d78feab9ced6c25735b3740a2309d96cb5d57fea729a9639d1},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{248, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h11974f58c95f8c44522f8359ae5e942577b8fb575a2ba18ff383df71, 224'h6c141327f9e405729c300f16b301de140c8df92c05637db952216e4c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{249, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009d5d514b884b4d892e92e373663e394901e483eca8c9bcd780910c82, 224'h7da1cd12c575744ff70cfb3513c5eabc0e3632cf2ce50ecf0f55c822},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{250, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f68c1b642a35a1988f6c2fa77a5533a2f635abf02c6748f5a2b9d1de, 224'h63ee52149fec97e52b2da4556fe28acf8f598636455f322cc9f47175},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{251, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h48948b8dd7e62760af368fdc3c225afdbfb6b98a1125d8aeb62419df, 232'h00bf889dd8eca1456c24d88abc16a5dc0217d3ac72b0e57935bb803550},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{252, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0d002750cc80c0f5a6b2b1e6e08afafb4840cbdef6e32b726a4c1959, 232'h00ee4095e31b594d159691777ff1f616989a65c4572b264215806f9268},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{253, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0977b6caba191d7cbe0b5319917f2748304e66577202335842e009cf, 232'h00b0680b5d606ef9baa292f6bffdc84c11c59299854b4624539c2efc74},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{254, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h023a1d2a8e49deac352acb3a6a758070b5c8a4e75fcbaffd9f32e862, 224'h5d2d511ed37cf7d023a5335c48fc2f63cf0733a1a786c49ae929ce5b},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{255, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c7cbad38e1c76603254dc2e9fd69332d0ef8f1a5879edb5be1bb578b, 232'h00dddcf1aa863f291c0a287fa1d0159dabfa7d98e646596e8ac41f1b66},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{256, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5c845a275521649bde9e3bfa07d6ca528f6e143d19e97b1e9e305e71, 224'h60b4bd522c44b4c32e87b11b6b80b2061da98b4cf5c56dbf5f0651dc},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{257, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h260418182c819de5bdb8851c5ac937ab8d83ab70640010f7eeae13f4, 224'h034c2f5ffaa2b4f1f111f4758e5adfbab5b7cfecfa48c8d88f5b6816},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{258, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0346d6521c74bfb34342c4b03c067d3cdfe35d3ea121580668301431, 224'h571dc84cc071e25b98d47c87edd3f6db73f995e5a4fa038760c43cc3},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{259, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f6d5049e2f0377f24fd3edd8ec14947251c9d687a4ec104f36b9238f, 224'h713a07b0dd9aa2b08c30d9167b0373b852595579a7dfc48199056178},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{260, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a7994553f1a793ebce2dfdcd357d3e4a01d0f7c1caaa9099fbb4b07a, 232'h00d8f771084d362ef2a0dee50496e450b6e812e40c2e6d342495571508},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{261, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h43236a22ba681bd71f99a8ee2b425b784ba6ff55cae154bf1b8ef454, 224'h09cffb77306a5ea7675578bcfa2d2142c9dbd84401e09f78ec29fa74},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{262, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008c63dae1f19d97135df18f8cf1a09e528b11ed2eac9f4b340621c73d, 224'h3095be2232fe57d372796cc0c846445836ff35f25a38ce13585858b2},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{263, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008005bcb6b955f80b2a2b6e45d86154c561b543083ab065b50bffb499, 232'h00e6515a9eb3fd8138ca117515d0f9a6549f226a72cccd49741adffec1},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{264, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00be66cc8eb0d9e5dd7ef6c754018502e7371c0b0db97cce378b9aa355, 224'h562b771c5104385878c3b918379b101ac888b1f15f0f52d15e0a92ba},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{265, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f42940ed7287b281f00c795abd671feffded542fc63c4ecfc7336427, 232'h009049e62c464723f50c265fdbcf7c6794b5294a58b3100e82ad9cd724},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{266, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d0b092867808c7d3b34fec07c4ebe8324a1a4ff2bfc2e20aaffbd248, 224'h4eb922b3de3bd244938adb20e21cdd560030d13cc0191c37ccd38e28},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{267, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a73472e1f303bfe50128770c9134bd93af9b064f9b782a45dd85c33c, 232'h00da4b8bd6e2ba5c635dcaf9a7d2bf774b10c2b09ba074cdc58d9c8da2},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{268, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009832ae82080ec02833e3eae913f7a98eb9e2d05133e5f2c7fa20479d, 224'h0e90c676df7737adb84e54cda47af9f5d6ab2f34eaec837b628f646e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{269, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3eac05a747f43988dab987f487fbca8003e5c7e9bb580634afef6e03, 232'h00dd656679e1c1800f8a258781f45489e6630a6d934b3e2a05d41a0c4f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{270, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5f3a639c163daaf3e2c0d7d1a3ca82ebe42951491114b6e257e28f69, 232'h00ea0e12e23d485a932f1aee974761b0e0c9c3d5ba1822ab646819886a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{271, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c0ad06ec18c4ed4469c5f4f4be4bfb41b6fc024456b2eed1d8096a75, 224'h45e08a93ae4e33bdf35379161843266ecd2f200ce292ac99894748ef},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{272, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0f5a1bb9c572a6ddfe5072de6a077b1490096a88cb2be9af8d976483, 232'h0092e7258459df848ffbcc7fbfa99fdf4db16b734dc5b9701427034f80},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{273, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a097b8422452dcb2a93ae32ff8d6befc31d76051704b1023ac5c7645, 232'h00f4faaf5f0dc78023885823c5547a59320bed2eb2eb3b948d07ce49a9},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{274, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7b4d49838bffa979d0d9772f8af39340023a6b11a0e2173ce92d1b8e, 232'h00f878af3f516288abf324b0c52dbc2d7106d2dc397871374bd144c272},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{275, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00feda6c1c40c483f87f4586d23381a71a6b051ce28916f199295eaed3, 224'h75be57d1b46ff0364308db2725b19bcc1ce820cf57e37f825d30e199},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{276, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009969b8d03ed1313ecfd1739e4c9234c0e7287f15839ea1e6feed50b1, 224'h45f6a820ac45d835ecdd52c836f157ab2b9279a560d2fe966ee23a4e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{277, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a62e952192d3a9dbfc2ab20c57c719bf52eef859d994c860a9564f12, 232'h00be1007b52e9308bde867f380f0bd3002554d8ac854f9db3d4a7d6898},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{278, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f526b9288e25aaea8d657ec7a4ebde46d8adc4c6d909fcfd7e2dcdb0, 224'h5d10087d1263db5259579e9987b410001b774f81c3e489df85b2715e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{279, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c5ff7ab638b6702535ea719e7c2f7753c53c1611c5919868fb708b00, 232'h00ab29aac043d35847280a3d77590ae93a4b26db18238a53c67cbd162b},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{280, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e69b43a68f452d26516e1316d54cd51416a047d42945350cdc506518, 224'h66d1abd5aa58eccf9ebe9391cce8cefab162a9130439235f051fc437},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{281, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0c6822e256d0190b4962c5b4bfdabce10d277cd347caf0850892288f, 224'h3f59727e4d9e3b92f4b0ce710c5112caa18e4051cc71450f6989cb9a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{282, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00850b43461e107174a77a4f9a3011e03854d6b5b4a0a6250e2fc472a2, 224'h0e7da9a21a2373d0944031fd121dce0594aa8721da1269f846747f59},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{283, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a6e142069366be8c48a7b651ec45b0e2dd9d79701108c35997ca1a4b, 224'h20b576040b9f3e73ae7ff3af223e34df82dce8533bf1901486a8b3d2},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{284, 1'b1, 0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h58e4c5558f2d4d2baee361da0e907e068bbc697b3abdbae29474084e, 232'h00951de902c7af71b5d7a3c6117d258242a04a8661bfdd4d047694f7fa},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{285, 1'b1, 0, 232'h00d37fb4abe8c504504f010539eb764c10c14250645e846eaf41b99953, 232'h00c4e2c1c277056982c5b81305ed3110a064ff6ae8e0545f0c35ff8871, 120'h00e95c1f470fc1ec22d6baa3a3d5c1, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=120b(15B), s=232b(29B)
  '{286, 1'b0, 0, 232'h00d37fb4abe8c504504f010539eb764c10c14250645e846eaf41b99953, 232'h00c4e2c1c277056982c5b81305ed3110a064ff6ae8e0545f0c35ff8871, 232'h00fffffffffffffffffffffffffffffffefffffffffffffffffffffffe, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{287, 1'b1, 0, 232'h00d9aac11d0277a4b23514c4d02a483e922dc40c92a774b8c62179690b, 232'h009cfe0c9b060b1a49598318631668083e4cf34e4bab29d14d81c2b049, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3b},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{288, 1'b1, 0, 232'h00c359b31b3ee10cc0bab7d21f0cc5cecb632186e8ca608a74f921986f, 224'h27787cc204c5ed561897c14961f7827b5f97395996de6cff87862771, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{289, 1'b1, 0, 232'h00b21fde4e399d8cbf8cbb8ea8ac770eb97ff85b018683433982ca2b35, 224'h3e7b4325b4319bbd71fe9c3e49c4daec895501afceaa554040129b71, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 232'h00bf19ab4d3ebf5a1a49d765909308daa88c2b7be3969db552ea30562b},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{290, 1'b1, 0, 232'h00fc0341bdbbce3beee1be9f02e46148af9da53128e0e3c45af1abe4c7, 232'h0092acfd718352e7107fe08ea6a35d8badcf54f57065dc4e8c9f2705d2, 8'h03, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{291, 1'b1, 0, 224'h50b14256f6ea50d9843bd9e2b4c2d9daf75f76ac4e4e757c712b3053, 224'h594d68e1683ec977b2efcc8a7ba6c46a0e6a668a03f4f50a3e21e4ce, 8'h03, 8'h03},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{292, 1'b1, 0, 224'h7801e48011fce2685a2f563faab34fff728ebb6e92eb029fef124eb5, 232'h00a9be2c1b86e99e44ef60e6c02a04a16cbd968482ed2ec4c1463efeef, 8'h03, 8'h04},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{293, 1'b0, 0, 224'h7801e48011fce2685a2f563faab34fff728ebb6e92eb029fef124eb5, 232'h00a9be2c1b86e99e44ef60e6c02a04a16cbd968482ed2ec4c1463efeef, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a40, 8'h04},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{294, 1'b0, 0, 224'h6cce004abbcdccdb3fda691e70a71a4d8a920219af2a20880f59c53d, 232'h0086023ea85caa2bebffcb9f360082e6264466ea065afb07820dfb1a9a, 8'h03, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c6f00c4},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{295, 1'b1, 0, 224'h5d1b27dd47711d7fa90b2651e202c240cad281ed803e1a3236c789fa, 224'h0ea5420664e2a8bd9cea3740218e23735ee2715f8130beb437419539, 16'h0100, 232'h00c993264c993264c993264c99326411d2e55b3214a8d67528812a55ab},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{296, 1'b1, 0, 232'h00ddf53cec8d9c6062904d2a04f790f4596c67696dd4f5422a3cb84c9c, 232'h00af10f2d1eb0e0ff28fa8e40a91d8d4addb20c085d635158de1a67bdd, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=56b(7B), s=224b(28B)
  '{297, 1'b1, 0, 232'h00f43b4a87dc12c65bf27f4b8610486402327adc0133c1db8adf4e3f9b, 232'h00a61aadb4c58ac0b5518d1c2929068eaa0d6a5d5f84dacf66e5b276ff, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{298, 1'b1, 0, 224'h6bd0a5dc98a6761a24d4e5e6c31187af8c7ed874d42af841806583b6, 224'h022e6bf9480c23d1be341f59b043afdaa76bad8622204fa84e26dd3e, 16'h0100, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{299, 1'b1, 0, 224'h75b65cd61449faf0d4bb2d2300b134757b714fbc4efbd6631e664cbf, 232'h00b488633f42e50b11c301bf3736a461286eccad2447180835d508deb2, 104'h062522bbd3ecbe7c39e93e7c24, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=104b(13B), s=232b(29B)
  '{300, 1'b1, 0, 232'h00bd18c7797449c64e9fc1ad2ca9c49132fc34b4741831fdbc6cbd87cf, 232'h00f830c108fd501bf9b7b3b898072397b9a6e72216db784c877882c87b, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c29bd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{301, 1'b1, 0, 232'h00af736667b618cfa5526f073f7048d5e6b672a05569cd2912bce8914d, 224'h6a030aa73fd79517ee8175800484f2dcebf02871825cc67c41b1a8fc, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{302, 1'b0, 0, 232'h00af736667b618cfa5526f073f7048d5e6b672a05569cd2912bce8914d, 224'h6a030aa73fd79517ee8175800484f2dcebf02871825cc67c41b1a8fc, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{303, 1'b0, 0, 232'h00aa2f981add5480e7f2a8ae50fc52258612ad6420a1a2cc2c252c1693, 224'h32c1ff19c331d3e52a98add7e7f4f8ac122ca961b8cbe4260ed83e4c, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{304, 1'b1, 0, 232'h008feb4b153b7dfe4081069ec708fdb161716ec3ed17c81efb1bb3e396, 232'h00bbc90cfae2c3957f2cec75239445239a1c0e9e0a032385d063f1d2ff, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{305, 1'b1, 0, 232'h00af2a29d356133f4d726c64e8ff7d80851649cf3e35d2b9de2725bbab, 224'h6d2199d9f3e0f0863e671deb987afdb25b6e6b7744bc53faa15cac53, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{306, 1'b1, 0, 224'h7bb0bc9529b06a424e8efbaafdec5aa339de5599f82ec9e195f0cede, 224'h381dc950caa8b0454fab70c57e06a15bc771b693ebb4013bc85b56ac, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{307, 1'b1, 0, 224'h2da3ea3145a1e68772e139f1b5d9b85e201de7df4775d5c4f7782596, 224'h4d3a2380099d7f3cf3ad18c1fb13ab1e054c097633fd51e67c1a9ca0, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00f18810142537c3fe231c073be9d0ee37a8010e002ba6f19e372a3f86},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{308, 1'b1, 0, 232'h00ffd40a19c09ce0a21124f163c72558e1f15a11aecde9dde08c465bce, 232'h00e3cc54426c7850ae17670e1cc19931e9d934610f42f456b8472a8047, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{309, 1'b1, 0, 224'h06081ee7d06ae8d4b84075e53264125b0efa082dc6e1d9190e9cd8f6, 224'h361012db570e279336fbc8f748d7d1c77967cc0ae188aedf8cb4d0f6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaa0f17407b4ad40d3e1b8392e81c29},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{310, 1'b1, 0, 232'h00f480a474e28f987e1e76e73c7a9c5c12307f5bdc99d97e515e71ae42, 224'h0e310ab3403eb44f8f17e217914d136c8e2341f71177052d4f07dcb3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h04d2a54e9e42beab49a152ec0764b823bd92a0bf4d6767e261bb4e3d},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{311, 1'b1, 0, 224'h4655a8b7d46613d3d8ace597a9d381b7d2e30c57aad490e413481105, 224'h4aca5463f0377db9c9638d280129cf14f5e60c8ebcef4c8ebdc9b15d, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00f9f9e7f101b4ea468eb78fd9ba89156454b414fc17d02840ca81ca78},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{312, 1'b1, 0, 224'h6c3c1069fb76da43e5a9ae1a69fb679740171f2b457956b13f5829c0, 224'h4f0b1000d41a56d96eca18a626d0636f20cee184f3d2f5b87ab68c4a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00be7ed7384bc8b90113e58ca87a68a06fc2fe5efa96f0a956733dc65c},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{313, 1'b1, 0, 232'h009a24375b03b78c20230867b842c680bdb88604fa93f7c59317348310, 224'h60090ff5dec7b6fb6df459befdfc5e9d440198e8610a267daa9548fa, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h79823515d525dc02f18810142537553a6da56048fb999d3fdff85f70},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{314, 1'b1, 0, 224'h71f01e6070a5bd694092417f75b1f1b35457421e9997fa5086dfef4b, 224'h2b8f67510ac820380907503b3bcdb89fdb5f2688434dba79d3a40a11, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h23515d525dc02f18810142537c3fc1ffd9a43852c262974a2a1640c8},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 0, 224'h453355214278474735b32b1d45c9a203421578c10acd426e9a569d5f, 224'h6b5655138346d0bef9cde0ebb97b4938e3c28dc612b4eaaba862182d, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h46a2baa4bb805e31020284a6f87f83ffb34870a584c52e94542c8190},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{316, 1'b1, 0, 232'h00fa86cdd0976acf06b0a7a3dcae70f287e62950d8874b32abcd59f755, 232'h00bd00817cea3c6b5e8d3266bef1f3df944fc4953e7a960902901ff380, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d525dc02f18810142537c3fe231b44eeebc76f3ab76829dc0fb7e7ff},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{317, 1'b1, 0, 224'h6fc6ce348cb17cf57fe18e21ed13e8f33e5a724bf87f151ea7579633, 232'h00bdd1fb53ba4ec9a477a6f3e5193003aaf462c857bc4a20bb62446552, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7d96ad58b0dea0aa5b2f5689fc4d2f3f919327bf633ae0b17d506e00},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{318, 1'b1, 0, 232'h0098f2f5da454958c7b04ef2220d45ed857a157d3874d033a25af6db87, 232'h0090c711d7574128fb7de7f316f7896b898670c97798d05a97f9eab7b0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00fb2d5ab161bd4154b65ead13f89a5e7f23264f7ec675c162faa0dc00},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{319, 1'b1, 0, 224'h3ccb08210d0b2283f3ccb779079bb160cee3cec9263d356565f770b3, 232'h009fb0edb83cae0b730fddd5c0d63e10a99e527497a58c18b84dae8e8e, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h78c4080a129be1ff118e039df4e8771bd400870015d378cf1b951fc3},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{320, 1'b1, 0, 224'h2dd3cd29db7616a6dc77bb1a66e849133b1408c540ee2ebb01e07bc4, 232'h00d3e5786401c4533e15697c6bf86e14def5088590c19aec9d96f8538a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h5f3f6b9c25e45c8089f2c6543d345037e17f2f7d4b7854ab399ee32e},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{321, 1'b1, 0, 224'h53e89d29406622bbaa1bcf7c980d523209646cc20a4b3104aa344264, 224'h7781d3de43413dfa061aa9b2d7c29eca9c8ed42b285fbcbbe016cc1e, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{322, 1'b1, 0, 224'h049c4d998c0f368ebf1a69274fddf807dae245b4d3144d696d813ed9, 232'h00a5d3f586315ee7f5b263efe47a1b0a2e94847242710370d92ceb24a4, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00855f5b2dc8e46ec428a593f73219cf65dae793e8346e30cc3701309c},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{323, 1'b1, 0, 224'h4b1b3c491443d1a45cbe5fb2f6ed36ac3ebde2a2456a7f9afe628dd7, 232'h00d328db165ee1110765797569b30b041984790ea3aa65bd0ba3341818, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{324, 1'b1, 0, 232'h00b19e1369acb5fc913d1ac6e92ee3770590c5a45ce52fdf64a9f651be, 224'h2fac7a017a6b6cfc1c381c9254564c1b929b3c101f89195a6d27907e, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0084a6c7513e5f48c07fffffffffff8713f3cba1293e4f3e95597fe6bd},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{325, 1'b1, 0, 232'h00d0c80d942da3dbe662467e1bcc69ceb322dc311152bf15557ed3f7af, 232'h00f7b627b0ba59524170527cc1161abdfa4a4a25dfd09c59a98db7ea04, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 0, 232'h00a781c88681c98aadf31e26541b9ab6efa52a49412cf7282944f13720, 232'h00b68ddeaf8a09af0b372b007e122d402e724fdcea1c619a80b32bfe5b, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d8ea27cbe9180fffffffffffffff3a43fa3662a899627950d4eb64bc},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{327, 1'b1, 0, 232'h00931606b9f180d16409efebc996bb1df442b84e19bcc9bed0e236cb64, 224'h50edd2162625a979a25b231fba17878b756a77c167223886613afb03, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{328, 1'b1, 0, 224'h1df7985b13decb2aa170b325ed2421d8d42474152b1040724ed7f28d, 224'h77ab5d47a2fb85754a3515682f20b3a47d13b26bd59b72f3bda83532, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00bfffffffffffffffffffffffffff3d87bb44c833bb384d0f224ccdde},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{329, 1'b1, 0, 232'h008a46670a9c9d3cf03a9e9d48525c75e572680a26278adc0888d5030f, 232'h008c88e59829d5a802c0245aa8b5641779877c5647ad2b9b2a736535eb, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{330, 1'b1, 0, 224'h16428097e6eb65688905678aae661f3d83b7e5ecc7787ed22fc029e8, 224'h68d62cb89be54d10ca5b575aa86f9c8fb475c6d90f59d4477595c01c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{331, 1'b1, 0, 224'h3fa563f806be913b57347adf8b1e862b7e0253bea701f6b201e57dca, 224'h0231cd68a2c24493deced00771e100bd001bc79902756d56d6ff87f1, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0096dafb0d7540b93b5790327082635cd8895e1e799d5d19f92b594056},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{332, 1'b1, 0, 232'h00feba9230660ac3fd64ae02f7306297aa4975436c0ad1105854e4066b, 232'h00ddcdba26679436b4e13f95d8f4f659142e7bf405c772e21788047b08, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h141a6efb8f6e19016b61c76573c9759309a18c16e48c136dca552602},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{333, 1'b0, 0, 232'h00feba9230660ac3fd64ae02f7306297aa4975436c0ad1105854e4066b, 224'h223245d9986bc94b1ec06a270b09a6ead1840bfa388d1de877fb84f9, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h141a6efb8f6e19016b61c76573c9759309a18c16e48c136dca552602},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{334, 1'b0, 0, 216'h25094ea9e4ce76d8c47356e4ae604eb6469669b0161fff805a765f, 224'h6f807430f186ba63ffa0f315be721ec43baef24b8fba10b04f19189f, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=0b(0B), x=216b(27B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{335, 1'b1, 0, 224'h754267d9f090524d4c97bb1a5622e0c9f804dfd70cc68d9872f0a4f8, 224'h708c24a49b81307db458c020fc7374770858faaea1d6ee37bf7beae3, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{336, 1'b1, 0, 224'h75a0d5291f48c17b4029baaea4d5796bda7c9d5802d534c0c265794a, 232'h00c93769dcaf7965f3c12864f50ccb22f10f193d5f0f7c33449131d2c4, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{337, 1'b1, 0, 232'h00d357674da166e0f4a058203df23b8f8ada82858034355d23aff5a812, 232'h00edf6d5265ed40b6da2adbe9f8cb6050ebf61ebc0e56a10a1d6cf6e2e, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{338, 1'b1, 0, 232'h0085675f96009ddf740108f5bdb82523d59414d39b74e11570a6d0faa3, 224'h13cd5841a8e2a3e3ebd099b43205ca46664a6e6cf19481e8552fb4d8, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{339, 1'b1, 0, 232'h00c1678bddce5f00e4f41ebcab86f801b4dc050a1b2da8f9747b5abfc9, 232'h00f1cf0d67d9c93456988a004dbcb8e95d17dde4070577e51d881d8859, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 0, 224'h09d2cfd575986bfe1a7420c7dabc0476e0dd13e54e01aa6f97b9e027, 224'h464ba5b84c4d92ed9fddd0bbcb2382f0e9b9d5bb201b2ea8eb8d3a50, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{341, 1'b1, 0, 216'h6fcc244352869febdc7425204f7b297ca85d5b0da8aa6ffe871980, 224'h62feef58d8c5a878d0255cd547af4f132906555017c330648d5b1ae4, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=0b(0B), x=216b(27B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{342, 1'b1, 0, 224'h0171e08f58fbf9812ae32570c2102e843968f5f35c596ff8591b03a6, 224'h6c07f75d9ecc5e39dda090ae92157e5d86fcf1a8c395490a446dc7ff, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{343, 1'b1, 0, 224'h330586236257b3dabb8fa249fc6a65fe0f97e4d51c162028e535b74d, 224'h20101ba5cc9967511f794fa7c7f6114d40e14b7dc589148bdb1c275a, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{344, 1'b1, 0, 232'h008044b73305e9f59021dbd0ce462d0d8a9b22e75887c56505c9c94c2e, 224'h6291a5c5364bad138d3ac3b538f77b266903bf71b6d4cc25ac0b6f12, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{345, 1'b1, 0, 224'h6fdbd44d22532a8803568b512f27c107572a4f0e99c90ab15d6c1bc7, 224'h014e5943da516a92cf6cf1ffb4f859bc93e5a8dd9f9b1906d69acd92, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{346, 1'b1, 0, 224'h1b9a838b8899a5c7b9d982bcc080787521d8334fdbd2bb544ab10f46, 224'h76548c21fd012875c5364e1552a03a1ea237a2f1adafe6279419877d, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=0b(0B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{347, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{348, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 232'h00f18810142537c3fe231c073be9d0ee37a8010e002ba6f19e372a3f86, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{349, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{350, 1'b0, 0, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 232'h00f18810142537c3fe231c073be9d0ee37a8010e002ba6f19e372a3f86, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{351, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h474b086cf4754c270d20f88be569b7d7b6eb6e55de6ce21382160e81, 224'h60692fdb35b4cb824a2729fb175f709d06bc9f4e8bbb4b1058c53788},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{352, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00dde359fe51a6d8ca9aec41e3376bd3e9fff8a41a3e44a64db81d6326, 232'h00a1c29d577309f7135b688b1990433fb45c5dc17a021557272c1256fc},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{353, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h0cdc4a54a091e61e0f764ddb12ffb243f457ad571a8ae7999caa0f06, 232'h00d5cdd524f2092bcbe2fc7c328b0876d436d9190058700af370dab0b7},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{354, 1'b1, 0, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h6efa32457e09b8abe22168501bc4ae051d2294674114a9dca94c51ae, 224'h3173b652c78324b877dc5bdfe80324aeb01b171fd2626124a44f0b36},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{355, 1'b1, 0, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h41a3e0370cf8148bccbdd03a7e763d382695263da11b9470b0e103d6, 232'h0087a612990d0a4a9f811e20ac520a3476d91848444cccc4c8138ad5d6},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{356, 1'b1, 0, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h6f138512bf05addbb536b976b9125e1228f43f32f766325d1c270e16, 224'h556205464ff65c9a5d4d9475167059863835644b06862f1b49cca20c},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{357, 1'b1, 0, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h00840dccce1760f476240b516d5cfbf9a10fbd44b25c68fd69a96f67a3, 232'h00b79884b6495a1c65f07853fc5d56ac06b84366bddb3ddf56b0fc9328},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{358, 1'b1, 0, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00949e76e0e35be5a08fcb60d8f86ecb0c650fc9b37ecd61a059649315, 232'h00cd870903fc1437d59e43eade139aa8eb717039d2e8d3282f27d484f0},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{359, 1'b1, 0, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00a6364e1e4dd41327b4f88a9998412bf168551acc561357d2bbfd2aaf, 232'h00f5e48ced76655eb729f4371d20f5d4ec53a23844313423063bb85fba},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{360, 1'b1, 0, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00f572bd069ffef726222db033664205220bf694f374282c795959945f, 232'h00ca942ef4fd6becd3bc4c3280ca29b84c8d29555dda402a50af1d7665},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{361, 1'b1, 0, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00e8b29401b22688776f8b24951f239893e12d822868dbbe1f6bc860ee, 232'h00bfefb3641875aa10c3e8468665071658d0ab312cdf8f9a669bd82a7a},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{362, 1'b1, 0, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h291d8cc81f715fd52a74168946ed2bf2d692dae0955249e4cdad3209, 232'h00ef56a69ebd78125a4ca12bdacd193e2111a35158d5d78b5d30460a34},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{363, 1'b1, 0, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00f5123a9f9212f64b8c607cfd5b0418f3694ce5ef4d161186afac7d30, 224'h44c4b5d7647dfc1ed10f1d8d9283d4bca6961a4ea78cf1cad632f95b},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{364, 1'b1, 0, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h6119c72d6d5fe72d181614d3d40b36eec756ca7d9e4f2ab3095d52a4, 232'h00fbbaf5bb4a97b6096792f17f95b116a645fe1c62fa1d83e969c0e8d6},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{365, 1'b1, 0, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 232'h008c3d675a759d30b8afcbee3f37746c226eb992177f8d76f162d4093e, 224'h643322d3f37ba532e7e5f0f0c14b691a3678075c03281203eb529745},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{366, 1'b1, 0, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 232'h00e1f7acc96fd3eafc29991165223b0b899c2b04cc239372eef4d060a5, 224'h2a0b6f214fa197cfbe834a4f80a74de9748e62f2a894214fe92bdeeb},  // lens: hash=0b(0B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{367, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00ab49a92649a5b95bee1a0e4dd897d5f5aae7581faa41673ad4d18eb6, 224'h5df9e1a65ad72a88f58b0b711e162c6de169ade7106c01571486c7df},  // lens: hash=0b(0B), x=224b(28B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{368, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00b3edcc316dd5cbe6cd0054e48bc1a77e55cc4cf3dddbf552ffc4e929, 232'h00cf4de654980e88f7908109c5f637113cb03bdf8ba5443dda852e6313},  // lens: hash=0b(0B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{369, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h32538b93b71e7ea2b3cef6027271e0037b84f3818a0727accaaea6d9, 232'h00e6225061a7d76b93c6562de31d50608444a533bb5853b8ab94160fea},  // lens: hash=0b(0B), x=224b(28B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{370, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 232'h00846e6b4ae059cf673ac2f424c07be6b64456554effd14d4a0a85d5d1, 232'h00c67353e85fdfb421fb3abb014f1d3d21a8b744ba146e4709e722a5e6},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{371, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 232'h0095073bb824196016092413631dd4208a571744d0030dd54352611921, 224'h100ef7ac960937e740f868bf9b37c6845317ab1865ce13881ce5156b},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{372, 1'b1, 0, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h3186a92aa760960996aea13f3137acf00b82b2b2036e607ec9c44b67, 224'h1835944e96b6ca1f445cf3350f105a97a37252f85cf6d8e628c96a02},  // lens: hash=0b(0B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{373, 1'b1, 0, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00cdb43f063ed3ce20f94e453d40e9d7de39936906484114c307078e22, 224'h26d2436f2f66a954010e580b95e21a174a4b667aa8249f2676fe1be7},  // lens: hash=0b(0B), x=200b(25B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{374, 1'b1, 0, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00b29a2bfe9fab394b34550483f3cc811d9b86345f6f8e35d6a6bb0b34, 224'h26120ea06b1910c44bc370cd0479c6addc5bce896c4a606810194e2e},  // lens: hash=0b(0B), x=200b(25B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{375, 1'b1, 0, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00ac247dff26016109d28200505270cf2d2c2b06067bd5d330a1c2a41a, 232'h00910a8d69da5d6a508c88aad4f091ed5b5286d029c1095fc57af2a106},  // lens: hash=0b(0B), x=200b(25B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{376, 1'b1, 0, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h00bfdbfcd3bee9803c5060dbc69d6749fb5e4dc40a1c00002e0d235354, 232'h00a84a6ff4c2ef80c074c8a8a9305e79e0e75321b9afab9348c02a7e29},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{377, 1'b1, 0, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h20fd72eb73edda9cb0aca2473c5c582c78318b0705a9a6d7180ac767, 232'h00b07a3e773fa28f513202b69903b5cc65f2b4f7714b5b28c83b52bedd},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{378, 1'b1, 0, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h0086aa1eba72a1aca7dd83cb2c2659241d12fd8ac17cbd798cc44afabb, 224'h66e0a66a78c6c31ce99e45162a0b4757deff5ed80be8348283f1b7a5},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{379, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h01cfaa7ccae0522b5363b48ab1fa5e0e102666f2ac5218c5b32523d3, 232'h00a61491de2a4a05bda0bf2769453faa845451207c4dd3a95aab169b0c},  // lens: hash=0b(0B), x=232b(29B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{380, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h500c9d08a0ab52d35fe5cf9d4eddea0eb8cc00e8e8db0a29a512de10, 224'h482d0f78f2808e83f10bee9fad61f4bdba83ab9a4f7d71c9b7083e13},  // lens: hash=0b(0B), x=232b(29B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{381, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h75bf80b060ff123c0e525c98ca74fa82d716a09c21d67accd34a60bc, 232'h00eda7a9644563a349ff3a2483b6e7563f0aa4c4d319551ca0c3bd1fe4},  // lens: hash=0b(0B), x=232b(29B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{382, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h3ef832679f6277b901b6a986833d03e4b574d23fd73edfd936689761, 232'h00e82af05ebafe22ccd384336c9530738036d99f17b62ef3dfc4e0948b},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{383, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h009504b624b116a2c28efa037e35581c71b2e7d01f30d8f68946c13e88, 232'h008082639374a8d5e067a6df09d6df11a972967a081a5307a3b7f1785b},  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{384, 1'b1, 0, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h2eb5db8a9e1c82ed4ce643c953c9f11c3de264ef92d7607c91dbce76, 232'h00b6a97c943aa7a62b5783786356f7b75b36b88356eb62d5a3d15a7029}  // lens: hash=0b(0B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
};
`endif
