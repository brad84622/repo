`ifndef WYCHERPROOF_SECP256R1_SHA3512_SV
`define WYCHERPROOF_SECP256R1_SHA3512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp256r1_sha3512;

localparam int TEST_VECTORS_SECP256R1_SHA3512_NUM = 99;

ecdsa_vector_secp256r1_sha3512 test_vectors_secp256r1_sha3512 [] = '{
  '{144, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{230, 1'b1, 512'h940016e8f13841a9f29c65adbe20d7c6ac3d2a8817aa34e44be00ccc67db4f935bab243b106b6f3d68b875b328a96379ad7491c16643ef7d37225aaabc79bfb8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h64a1aab5000d0e804f3e2fc02bdee9be8ff312334e2ba16d11547c97711c898e, 256'h3d4e6c69176bb9e30eec304a30d982cb3f6073a2273f36b67b1b284899b08163},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{240, 1'b1, 512'hb1fe8fe86f9994808c00000000f313a999ae7b5281bcacf933f05e4c8d526e761afa3141e9efefe959438620220c28bbad7047a6c1a98f95520baeb1d7af6278, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h33b2abf92021a14fd1e5293008c8aff551fd4a0cacaf8ec6e147f40d0f521cb0, 256'h4d0d3ed085477a4dc7fd86d242905637a71700ffd4c22cf962a67e9ae32b8877},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{241, 1'b1, 512'hfa3ef856182ec646db7300000000241a0e98fb88ce661de43bfd86f1c929391ee9ce6c05612b1609d6b8466a9c4d0af24ccb440f463cd18addf4674adb2f94ea, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h717f5185242ac57215d8713f902cf9012f45dba76b8e7e51c67b71e6de10f0d8, 256'h28a9ad765a6b1248807be126b9eee01e8e2d65d8528cb28f0d45763f507d97f0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{242, 1'b1, 512'hed19e69c6f4de76b35ce6c00000000ad94175b8ad5f1fb69995d7d87abd893772b81ff83fd6caa25d1fe69b0317ec4068cdddac49512e6bf12d9cd8ce9a951c7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4e57dbece14d3d279f1e831777b28401d2990c4ae477eebb997b583e82f29c54, 256'h3e41fe090c8f14b8af7fd39c2628869258cf05b0e289b6692602c10cdcc8dd83},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{244, 1'b1, 512'ha8f658c6632e4f474a6f1af1b9000000000048ac2a6121c8add714fb8cce854dbf1871b07a75008a42baa6cef01b4875eba4bc9327b41503cb36ac20f9354238, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1c66a303f7f548ff4c17ce6c6038879cb9d47abbb71ad69a798d0d8a99518dcd, 256'h485ee205c6fa3ffe5411948dff2351ab9bbbc20ca419d6182da77f5579058749},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{246, 1'b1, 512'h9490ebaece67e31eca85b20871120000000077b2785e29958e0ab90faf8fcca953b142d51892ae5362246dc07a066ff6a4c9fed90a79fb59abdb7c8a888a9652, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h67afdc527b0003c8400ade54df5663635f811950cb34ea77435c0ce400365249, 256'h7afa3d39b8a7e52ce768e466db6da41a354c12ea2f677bf05a24fc689e347323},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{253, 1'b1, 512'h7da7793b2bed3ce23ef7f1c04376791fa03f741f650000000008744fe10ac37fab4edf76492a339fe79e56ef75aee6c3169a0a61e3cb27e74666a4fe4184526c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h257e760a54637387b443f829f1a5802c7fc92bdf033039acf68e1acea0cbcdbe, 256'h25087f120467a80cc07efb7bb27ae68d8569a38fe2908282c3c7a310322761c5},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{254, 1'b1, 512'h48cd33f55583315ab2131d5db1f9cfcb0590b13a266700000000c9bd5d6fbcdf457e3bffd7b4875145a47be68b99a201b93b8685e80d61ce692a913be1183569, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1869c821e271838453c88c4a867df2301d27662b72d9385bacb6740ab6d6b5c3, 256'h22ccc9a0493116556d9ffc7582253c581452d717a7e00618dce21f46f5b64fd0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{261, 1'b1, 512'h57003aeb6ad8b84b54cdddb9243c65d8fd07ad1ffdd35f11c319f06394000000000aa9393490e8dcaf1c1e53ab5a7b2dfc0bd1dff4d0fc1e0c9dd5cbb035748e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h457ff86369e4efd69592b161aea2b09153f37cf69006907a7558998ab34b38a4, 256'h12692ffc569849dc8e3b9fd2cd7c6f42207bb4c07832d490c9d35a702665ce58},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{263, 1'b1, 512'hdfe80a6b887fa09cbdc8bb94300a4ad38f0380331a18c0a0b62708e590dd3800000000d364091041bb72f35391e792802f5c23fd676d0775e56ac2e41880d92d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h59baaba3992dab0b594a2e9fbc4c344cfdabe7868e4e77f47a310d94916d30ce, 256'h20b16c383085ee74402157d4f2da5f7e3e995dbbf53ee50985d4f7096882edda},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{265, 1'b1, 512'h519e4709f22b7ec44e321f4d403bdde7f532392786df003ecda243880f79f899f7000000000e3e6d749c0a602d959e0fd13a8a491554d233b9dcce6cac4ff3fa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6ac18c06081a51ac5fb6d0a0735af510dd0ad529206e7fc0c1b6d0ea36cec4a8, 256'h64d49524cc26ef8eda21ad5f2c371203d6eef8ddfa5da7a6c37d86f29efc1fca},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{267, 1'b1, 512'h2cd7eb20ee13fc351891dc4acccbc978161cc1b1e0cb95127485ff132176a972377cdb00000000add5eee3b407ef394da0255f21b9b8ca144d7e76fb075c6bc1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h455f1c4406b598fc828ddb3bc77df7ad04baad399fb4975f542b19aeedfd5a11, 256'h4e0555d9bf4211d3ab173e2e6c7edb990867f8f982f6afc1b4b6732ee96a0af0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{273, 1'b1, 512'h4025a46ad55fab109832d892d397d6e50c9c0aaf7136c275c259a6a61333a7e139b394a288148e32c200000000a3d26314f0694c5db5058ee34dfdd8fc2af9f2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7973333617680ff89798c6b64bb42f436be7771887c2d14a98dd3397e6896e0a, 256'h11b70b23a62fd9ce1b27c1b669c851187c09e9081f0aa6ae011411425f694929},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{276, 1'b1, 512'he68fbb72e90ec509836476f39f26d3f65c5deffafd5b86448457438ee0c621fc8f97e83c77ecd131ff1e33e6000000007c2a942574c7da923726d5304e0de79f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h51adf43cda1a938e1deb5fe08ab28df1e607f25fb2e98913d2579420b63056e6, 256'h3b8920181a8ab6f9ea0a1814171db3eb4ff3d5fd9cbd2d9c1ec4018a7625562e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{278, 1'b1, 512'h1c0e382d29f7ce824206c57f19794f9e8abe01e6af45a57dc9c01184c7b956aba27c6536c48c0951e2540bf566ac000000006db962ed4d45bf0d0c1c6c806b4c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4b2e5a797d240cd8c80b424a41dc47eaad249fc642e3c5b4bc68328fc1e26fc5, 256'h117910985597a6f7482bec7632e94676c432684f16f7f3d09a90ff4ed6ad36db},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{279, 1'b1, 512'h92cc3187d3326341d51f43165add210d496557c7a27669692c21c2912bc85d13d22a15ce9f2dc8052f89cdb3444fb400000000da250c8d1d81c198686e0c62d4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h42bf9a164723ef3f5cb59b528966ae648e80291785a4e0067283a7af59795bb7, 256'h017e1d24962a34d850d94187d269836ad437396a0ff134067b1baedef69b5951},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{281, 1'b1, 512'h290ba1c9dd4ce7537613a8092317a721e35cf33f17d8c82bc20a765683871857d7a7f0f72e659928158b11760b339f16fa0000000065c91469026a04f6e368f6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h183c81ab34a7d7c6742ede4198f5c75ed7fb79e8315899ef0dd26f95e3c4ba26, 256'h73f0196e459eb980b6e7ac44d868ab632d6421d1788b9f9651fb827b1a8e5dcc},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{283, 1'b1, 512'h1827524c50d2a178cca81cdd33a0be182f764450e04af569ce80811e55ddf11bf9b04675631ccc24d816b26e407df93f288bae0000000040fb10fffd72f8f6b7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7c18891499af92cfa1db5538c7afbd44605b17dd0ede573206db85af23d3fe9d, 256'h28ceff96833996ebababef332b05372209844ddcc4c2134fd9311397e733b10a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{285, 1'b1, 512'haec77ef7d501e59ceb458f4b03194d730583d8282b6bb01ce0b0417143ca15c2059e8290afa26d6c1e38502d0b895bb4cb182dd4cb0000000097ca7caccc470f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4fb615772d56b6d1ba60f371eb04c557e0c9414c4eec00819c7647d91e7dee01, 256'h2623c6c4a3bffc596cb5f2f70a5a381942d350df04c35978f6607ddf7d57e4e3},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{287, 1'b1, 512'he1942b44674c9c247d1f5857111e24baa87afe02ae74ac9d1ac122c10ced967b6243fd3055a4de1d50b98e24831c9f613d767a3060f7f600000000e5461279bb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h08012cfd3713068d8ba6f3fa453be9da95afa6572a893882075ed5d64d62a417, 256'h3c5d1bf341823a4cca251cd67d43a6bcd6b5e47303082b7e54c80df5acbbac82},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{292, 1'b1, 512'he47ec71fc0cae21e08260f64fa9dc1a4c99ce92048144beeaf932a124c0f87a8b0db214e5424891f30a4cc0311efbb2d49807cc31733db9bd80f912800000000, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3b4c2fb773223c1dafa6d6de9ed2304dc25eea1fd487442a3a64ae8dc8f14927, 256'h56c21579e85fc9075c7601bd36ef8a3fa57d5bc7550c9a17bb8383e7fdbb366f},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{293, 1'b1, 512'hffffffff149aabbf287a78cde6477453f7f9c2310cd2d58ece43bb07019c69c965ca25e8df7696c97ee4ecd4966f7577eb41a60745d031a94f5856e1a5f95aa5, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h05276f6159e2853fc6884c2939997b5a3be7ae615dad7517d6006208111dd678, 256'h059ea3474bc6908c565dfb5bc72fd1a84231363cf78c4c317a061dbf1b03cc07},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{295, 1'b1, 512'h9481ffffffff6e35dfab283e61e8f9a49de1cda44cdf1e2680292ded627b16d9b566ac057cef4c3380ee126c020a6ae86ded132faef613440c54185ed5986dcd, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1c058daeb17f995cbaa4b02fc1ccf0a121fb7673d7b9b7bbaa2c9d850f9ba741, 256'h3e5400acc992698dbe9c41e25547c6ee08c841d6604de457558ee8af11d54446},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{296, 1'b1, 512'h2d8fbaffffffffb42e8498ddf2697ff4a2223fac0c486f05f57374d84dab9e8d13f52f6c898c8a7a74f2d48bee3cc16265e12a6dca3bee77c0ff0ee5e9af7e49, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7a6c6eb198bced25223fed630dbd2956c3799a21389e007efc23a0b3968f8aa5, 256'h4535354e8fb477d0be4a16f44719d94650ed4607eabe206848ba24322406c1d5},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{299, 1'b1, 512'h37837a8407b6fffffffffac5686980dc2ad1a556be4d1fcf5dc000a18139c2322fb6d35995be1b96f942fa8bcb31b6d4c0efcdb2febaad183b00f4967c63c04c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h480a6875b7bee4ed80f70206400df10264c38be42b07443c6ff19c0aab580444, 256'h78e3fa1c2fe11208c189a39e717b19a51f5172054891c083931861c7919d4745},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{308, 1'b1, 512'hdbab4c37e253fc1deaa9e71c035737ffffffff6e927ee1da438de0d1d5152cd6d0549d2b8172bfeb94749da7ff020aa760407bc5e12a5a099a45a301588b62c4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5e399962385aec963cb80dab6b5f5c341ce15e437142f4275ef9c210385348c1, 256'h18a8157a0976bb0e349a02134fad0d0286c40a5e43a47b49b5a03653e3ae9e19},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{313, 1'b1, 512'h55260440dd65e8c48db54c801af143d639f08a95ffffffff9f03419e88a5145c37a3193cc07c160404a9b7d489aa324965d89fc40fab65a71fae34c56afa395b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h25236b00a0a67e12ea781ae53a929e13c37994ddce784f3c0c33402a43b4a6f0, 256'h117331e5b39fe2a11f5c8bbfa5bb4fdc3659ac0a0efcd03a94362081a4c0e579},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{314, 1'b1, 512'h16438d031fffee5b56365cb1a8f4bc19eb046a111dffffffffc16998d3235c27ddbfe7f1e45105d70ecb963cf511b0e09daa505bc426260466ec6528fd48b88f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0f3564b771337bc8d494a04e4d0518f26d067d07c31689d5e27b503d3652117a, 256'h17144740db21874aa58c0de6a4cadb16c5d9230d4f4607980aabd161d21045ae},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{318, 1'b1, 512'hde8b1dea4af73e03d31712528653ece2fa048092693f2106acffffffffc4fbe785cc6cb125a5ca069dadd2dd809bc3c6246bc299c2bd84aaaef1085a561dd79a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3977465917472d3cb67d6fc8888834f26fa47c8d3a2c8e046f70680e3037a37e, 256'h785adced4f3d400b286ad7eb7bdf0b7c0f46d9e7268db5a34e740166caafd14a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{320, 1'b1, 512'h0a55bcbb94c925c397b334ec37bd5216789d87fc6589738cdccee4ffffffffbca7bb2e94ddb13839ef8da502b39ac80f25abca143e0add021592ea7a36ce83ff, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0162ba940a75c7a12574736d45d60bbb2c6ce7739b04429cc72352adea4666c3, 256'h4c686aaafb4f3615247ff06b97bd76d49b93f65b5f66c93fc2a8a22246536c24},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{323, 1'b1, 512'h9e670958749c5bbc0cacb1ee6c38e71eede821d75d84cc2fe1335af9f6ffffffff4e9613cec31f535c4c7bdab269d70a8d4b3bdffa3065d91435a4237cae96da, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0afdcdcf68669ecc53b019d7adbe8dc943f453b74451335a631a2a3dd5672f83, 256'h77ea833468953e14bd428663eebce4b3cdef41e9821704fb91d1515d20078e92},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{325, 1'b1, 512'h59f9626626a34d5491d567d0315894fb702c1d7a2ec677a2b595a772b20d8effffffff20557e965f33f606242a59aea4cd565aecb931664e51fee93a92ccaab6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4b3eeeaf50e9f9bae0bfe64e2776bf2db181ab44c763393136927827f3adb24e, 256'h317abec131eddf2117e27ea2bb4008e8fd0f4a32aa41f74eec7b1659c091fd9c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{327, 1'b1, 512'ha05bf269c6959e1000f754963c2ee746346fac0d57bb119d3cecfa3dfe702fef2cffffffffddcffafb72da48023b4eae3593eb7c3c2d758c1c6c5e4dc57d53bc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h270250c591cb20c7978d9f457104afa7c3484879cfdcf9dc6ac8e785e1fd20a0, 256'h09601dc597c123ed7e76bdbe2d146863bddcf357f9217713dfe1afd8f49891b6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{328, 1'b1, 512'h9695a59c40d735b329f1f9c2ffd974ea8e66af6c65a1f7242e1eb02ea6721f9460ffffffffff9327209276e0633e07c96c9a2950a09411d1eabeda48ba90c8c3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h729a17311a2fbf9f2325117b2cdac18fd6bbe3db4c5a1bd4e4f4f3d8f3d68dc7, 256'h48dd0269cb216e2792f3b410a781c9b10e59abdc553aae2a00d4038f44a2849e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{332, 1'b1, 512'h125406f9b34e4f63c0a2288bf6166292074a0fed2b2c47822bb885520f2db3e2c58186b926ffffffffee3b259d2c85d9ab10b9f10f7f3cab27a8f528b4a82ad8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h381458d6c40c888bf90aef1428bc968caace553f94287e7adaa48943dc55315d, 256'h1e0e1f75489a451fc7cc4bca61a0a7330a5b4dc4283df68e21798996d8c69bd4},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{335, 1'b1, 512'h4e29d13bd24e9f13d5e31ac769469a23d44278a67b110f7bab6095667a3a5180bc8124849e31af47ffffffff94e438c9abcb1301833210026c068417d2da4b20, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h61746df1d5f3d30403f5281767cb6601172b26564e97c35d4c68fb7426db4ffd, 256'h7ca2b0a4fb0d58a119a8df391ad3f2de47cb3b1a8fdf04d6ec235f639fe44080},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{339, 1'b1, 512'hf9db531c8bd06c7272a9ae2de6b4cac8e0281438eac5689c7f763241db7b88b4a6c71d53a3d03222f6195dffffffff0b690ef5a310f733b13a1bda4fe964a38e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h130fc664eccece7b71a0a9cadc5369fb5bd54ccc53fd2c515e5ef232acd1b965, 256'h4372a69ef34ec2b296dbe94c5e8a8881645b9c0f6b6c4270c19b81493eb59421},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{340, 1'b1, 512'h273f59b9ed631e0fc10467687508d817c2229d48e45efa2a6783290c6ab048c048a882eef2730e7456b3d4b6ffffffff0369568d9ede46d524123c6cdf78afb6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7b675a89f3165e2ad1f3ac4950898d17e7cd869df4ef58aa54901d51193f91f3, 256'h3a7ea099d7c2909ff4a5c3c286d9f7739f38b7e44605ea3f515fde117a4519ec},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{341, 1'b1, 512'he6ded1492cb08b685e2c14f2f11d4bb2fe1601c47019cdd5bb3a42aadbb88f1335fe76ecf455cde30b30e18d35ffffffff921892b8870a2d1248dcd97ed5449f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h393a056a5ce76dc161daf1a6a77afb72cacb809d4173b9126e636a01cf7ccea1, 256'h0859e4195124e11e40db391a7bf04f3ecd7dffe2a5629aac9374468fe8f1701b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{342, 1'b1, 512'hef9ce8e0e84c667ba940ccb1d3317daddea8b9888a2ef5b718605aeff060c7140522f73cdb7670b0e055a2646509ffffffff81c895857965435d4c4421eaaee8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2d9738a6e36c24a5dcde61ff7fa5ecb1e96e0077a4a183e8953745cb9461e5fa, 256'h55abb27fad179d132830f7e5dff0d26a63f0141fe2288b9ff7943c3a482ac124},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{343, 1'b1, 512'h388b354799942c6595ba49bc6bf8e7ca5c06c6ae8015c0f58e69192d96cc60e30696c1284ba98c1b22c5c7f23bf8e0ffffffff15f579e355c7258262f0fdfdfb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h460f528bb6f8adb55626c5166c4572a93c3825dd1a695822a81c9e75e37fe8fd, 256'h0197c8b83193110f0426a417fae7ec3b99fc669371f1e7debbbd3850f6956c14},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{344, 1'b1, 512'hc6bf307fea8c2799ef482911ac86779072e5757f934a3671ad8c5a9e372bb2ec8d318ee3bd0cc4460f9050c937a3409cffffffff81c81c22e9468fd07ec09f55, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2d13939455192c22b1f18f7ca82ad4265ec2c4dbd124ae4a2b0017984512c9e9, 256'h3d9e4fac784be61e2decb75a1f6768af21873eb49881849b936036b19187a734},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{348, 1'b1, 512'h4f34828f9520f17da9e588884a26df5ab85e8456184bb19001abc926a180c32a112ba4164e81d69b8fdaaf3c60619a7d1a5840b6ffffffff8748db5ab09c4a64, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2b7d769ea682af0be42866cf3ad8865b12d4b37c3708fb2ad0dc5c87eda10154, 256'h11d8c48ba6c400f7950f9dfd9ea65617b3765db0e79778bb079fbd7db67b68f8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{350, 1'b1, 512'h6a763ddd1f348cae57162f918abd67d536a03431ed29721e179403366c3fe64f1083d4a64cb7a9fddc7c5a3487675be4078be3b484ffffffff2d5a70dd12c49f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h56a5c2c2e803e66c5751fe8fb348822609b167478cad4030e7bf6120fd535bb0, 256'h7b3fee66768794c0b362f2d40ad64fdf03e0fb0e8a47f2034167aae2ca383c0e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{351, 1'b1, 512'h0844602883dbcf60972c8b943b5ea020ccb0d19c82eb86cb18d4225a79f97279539214d6e3df6ba6af165c9cd95b8b67a36b39bbd101ffffffff5a9aa9794dd2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h71bc399e5643a1d8e2afc317e78a2c43d76b6d87f17a5809a7b6d19f922c2e62, 256'h057e7615a2c9033ef0d1a3d3020977002395e196d3b8206c9afecfb98abd52d8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{356, 1'b1, 512'h3db47a2cad8a1c43f31ee677cef231cda0f3853901676c1732771602ccdcc294a38fb8df77d5e6e5737d4c8e05953aeb81edb39a25931717b3c154ffffffff9d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4456d6792ff7e4d27517113f309177c26ef3bf6482e131d43f9d8b80e954d61e, 256'h4ffbcc50a7a69dfce92a47410f8574f7b0abfc8b4c7f74ac0dc1c1183d393482},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{363, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0c5baefb69764c3a55e9d3ef10a76f652ffa697794ab91169878116d058420e3, 264'h00ccd7b9153694151ee2d05048e40fe072d8e0f481af5d3d0a9e8cf39e1ef7e0bb, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h27b4577ca009376f71303fd5dd227dcef5deb773ad5f5a84360644669ca249a5},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{364, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1a4cb39a674bf0bec4be1a5b035ae18634f4b681a330c1f91b42366a0a7c7532, 256'h0b3f8018da54a8d0db30f7c2b3f04dc011a4a1c383221e52187632a565e5795c, 8'h05, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{365, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1cd72095fd856cf29fafb81c25f7ff24dee34eeaeacc0025d512091b1f1e822b, 256'h427eb3bbb915209e064bfbe1a1798ff6dac8d0add6d753bff4f128fee7e00f89, 8'h05, 8'h03},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{366, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h697cd5856c8c347fdfbca4c2cb2fc1be12f1611f190333b80a5cf4e0f7d48dab, 256'h5d08740936bbc46c90b1da916d5ef39c3d9fb9092f579a43d911472022a7fa90, 8'h05, 8'h05},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{367, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h69d31ff52dbc0935508755cd48cf3f30f0ea78fb670048983be0ebacf4de1076, 256'h773c9dce9aa24b783d8688d63547dc987d4650f20c1179e6ae5d4f14f6d55cc1, 8'h05, 8'h06},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{376, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00cfac11bd4b7aa0a29309767eddd337d302f1f42ccab215171f9622992a671e4a, 256'h1451102ad100a24e6fb5cb130c69de2a61fa50f2d07a099d73ae96f971593588, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{377, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00cfac11bd4b7aa0a29309767eddd337d302f1f42ccab215171f9622992a671e4a, 256'h1451102ad100a24e6fb5cb130c69de2a61fa50f2d07a099d73ae96f971593588, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{378, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00ca99e8cacb96b9b73a7ecf478617269f08971c307aba958692381696c244443b, 256'h5c5df1f740db3016b0ad298997131cea685b2ba405c3b0f722c6992bdaa6fd3a, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{379, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h3c31be015178a9c3d3cae9103bf25bc11a709316d06ab46c01f884a8eb33da2e, 264'h0091f32a1352712508642c4774ea67049175161cb2bafd5524b813274b140f8e99, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{380, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h355d9c3f97a282ac17f7bc98373f271d6a2bc02eb964f13c1e2d7debff4a02fd, 256'h63282e78fb9b88f81413bcf95f16982d9f50e7f94a5d28685b41da997201db5e, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{381, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1c959964cabaa5ce966b95acda1c5264847a780426c878d716d73ae6621d3084, 264'h00d3fedfc4f9c3b8cc8bc6539b821ad208ec08d5737aaaf1801d666ddc37e54faf, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{383, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00987a839ec570964d3a1bfc6a0334e7328c1624677c66b8fef3a5e64d1178ddae, 256'h5577dfcd0fe00da9e1d8bb8bbd952aaa5bc10ecb14cae4e3f5e28c506bbc3a21, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{386, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h36c6faa9f6dca42ea8b0e6d02d36c3941582749251bfa88c35fc8a8e9ad51cda, 264'h00c44ce5f20f36b4ae75cc7291678dbff188cf8c838b8963eeb8b78891795a7364, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h2a06d743967a1330ca91cc46c9394512cc85b4f1b9355eb7f4bbe53a32b76cf4},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{390, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b034897e2a74a787e008b14c62882eaee0e6e53a1c8a58f709a54432713c20fd, 256'h28e07de2ca64b5e215d25d0530d7807df11b98bb39c26a2405388ac0b163fafc, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5f025bc7c717fdb28319587bb1a10fcead32935ea552ae4fb0fe33cdca6473d1},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{395, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h3c0c4d0ad0848d1335b12a8919d32fafc5f2b0d5c2f3cf6494b06ba8eb17cb29, 264'h00dd7054095454fdb519279cde10259ec5d9e5e4b5a8c4daca649a150f2dbf21ac, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h21f862ec50ef64b3bfbe5d774e20cc838320437725338a3b32fefe3ff159dded},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{396, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6cf91440818ea262b9376e23f7b530b9e44edf5bc6db1a67dd60cc722975d623, 256'h17c19e7d6ebc0cbdc89388242d604ae94ac4ca179ef2cd8bf33fbf738afcb39b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h43f0c5d8a1dec9677f7cbaee9c419907064086ee4a67147665fdfc7fe2b3bbda},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{397, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1b5afcf39888d2da7215f36421a85c4217b0ac883bf5957c2d066efd8bc89f18, 264'h00d8fb3b6aca0b3577a883948e016905065a3fdc13d6f433172ee0f16784e52c78, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h65e928c4f2ce2e1b3f3b1865ea62658a8960ca656f9a9eb198fcfabfd40d99c7},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{399, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2a1571ed0ffe39574d030b406f638bf88eea5b4b50754e93431fe0172fdf2fbc, 264'h00bc77f601dc6dbc88cc2b560e8cca5e738f2c769810b2c8762dab917adfe24535, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffffaaaaaaaaffffffffffffffffe9a2538f37b28a2c513dee40fecbb71a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{402, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00d533c620a8fd3d5a8342caba89eadc25907d1e9b6fea48ee8f806aa772f0c80f, 256'h70e09c022fa1139da32a456ec024949824477bf0bdbf603e8faccd6b205d263c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h66755a00638cdaec1c732513ca0234ece52545dac11f816e818f725b4f60aaf2},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{403, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h0091014bea8705a022972e12b176c96e84c0b61c05eb1c6f8c5c1db731d54d67e2, 264'h009060ef6c764d8d47ed5ebf8f6c23835cb89f8b056cdf7e457f9273b6477ece33, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h55a00c9fcdaebb6032513ca0234ecfffe98ebe492fdf02e48ca48e982beb3669},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{407, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00aa9d33c76ccd011ba23047a420840374b4fa3be480c65263d543baf2ccc6141e, 256'h5ed3b42ad9527869fae92914b82b952d2c31c8fcc85b4c100983096694285766, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h266666663bbbbbbbe6666666666666665b37902e023fab7c8f055d86e5cc41f4},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{410, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h4b7b9990a6c2c5a810107c09ee09cf3388c1a6e82aaa44c378d9886e2508c2e0, 264'h00867e7632fcc312fcfdc01fb6a579ce6aa6285563b1adbb3272f0e122f9de73e3, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffff55555555ffffffffffffffffd344a71e6f651458a27bdc81fd976e37},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{411, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h568426540e19be6404e6cb4745fc7a943c0c059d7c7baf3bc4fc782e9aedf2de, 264'h00ba7fb20ad12a886c53945d3cdb019afa8b0d58ed307d55f556acf79ec89012d5, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h3fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192aa},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{412, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1bebc1a6823107d1263219e36d2ec1957d20b0b450b481c9de46ea9294d48b66, 256'h72b7a811af9528e61199f4a2a7f30d8685f5a04767b59276e65a732e8f3950a1, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5d8ecd64a4eeba466815ddf3a4de9a8e6abd9c5db0a01eb80343553da648428f},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{415, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h69aac6897b0457e54cac25f24590be255d352a20055004e7caa7cbb430b3c90f, 264'h009113bffe220db9143e38514da0481df67f1717c58aab1a189fb9d4f6e53c3900, 8'h01, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=256b(32B)
  '{417, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b282b1b5bc00c2bb18f28ce678e1cd48c8ced8335af5d8e4abd3d7a7d3616f56, 256'h3d47a55ddc11e966fde2bd87b028e62fc8133def824e3e00528f2442908fe84c, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{418, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00facbd6f5e996284a53cb1ca41ffc4eb0a3fd73b73c730194011169b9ada14519, 264'h00c5491ede60614d823b491198df7bc6c6768e064e0e43b7f053ab8f279cd4f4ec, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{421, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0754de71bd21f14f4927bdab77efc57f148b36275c305a86c1d7a0dcfd53bab4, 264'h00989fc99bc725da84197c2f284ecc6030489eda77ef92f8680130622b631af2b3, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{422, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h008aad84fd5d52afd531f1068fb7a10bb365faefa89975597187470d04a8c9c8b3, 256'h27258e32d19cd58ddfd35bd7ea1f063c77c61b7879451bdd3e8f44cbf40241a2, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{423, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b4a01ec7b10acff3dace05222fae05c75368a375d8ce1faf4a1b2def1ab715ab, 256'h61a6642e82ff950f373ace5c0cc298639ab9ae739e4614a93fb1122ee16d922f, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{424, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h4efc2bef42b11e0929edca3b025f01b1fa37aceef4cd3e8c2d4beab500856af8, 256'h7716828fc1788c881ae39f534c3e270ca869a578210b5dad8a8938691d0c4b73, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{427, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00efd3bd1299d4b2bb0afbce2afd90792d8c72e1d29c6092e4681540420664e275, 256'h390a4dbb20d10f7360c5b794564dcd443bb1df94bf6b1f4be5909a22a6a534ba, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{428, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00dae9cf165867da6482ede84bfc5b94375529bcb953f26d0cd68fc877088f78d9, 256'h51cadc9f61c55f8e2a04dbaae1251fd15cb12df9bcd072a51971127eaa6ce612, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{429, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h008418924e94161d350c9fe8dc1cc087de4b4491d0bc694a6862df4e8a555f9afb, 264'h00b0b391af97b0dacbdceb7a982781d0090978efbf76b8e6914250e92ade9a6126, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{430, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{432, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{435, 1'b1, 512'h86fe1b4ea7ac8e339d04e40087534c61e245dd4a0c22754a0622642bba56de900b2d431e859a36b1a5ff71aee560522eb0d3251e018c2cb6a10b82031cfd37f2, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h532d672c307da2891720d11422035ea25771f4fce0dc9948d754ca4f66ef36bb, 256'h4f296181799d3e6780086d6908ab8642711bd406e481b0ce3af1c44b9f098496},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{437, 1'b1, 512'h7d795fe6a97761d89b35f64e09555951f6ec2a669a9fa03481c100ae158f183e2171e142437d2c3a42352108a22a7e3d797beaf6c3075db419b6f4acca479c83, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h6637f14369d1dd112c5691969fcc867e64bafb1f5d8f917a9acf8ecf1dc95754, 256'h457b4a8bdd1c047b12826897991241700dad09666b4f410a56993023b098fd1e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{442, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h284fe5f1c86a55fcb3c27a12d82d794eab9a0d76d1fdc4f25df5a9bf52e8e768, 256'h7aaa75e5a7948be66f06ce52fc3e4916fc93514b08c51f84b73839d2c05acf58},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{447, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'h670ce60d0fc7224c8d06f3b01c4416ee0b3ac12f0cff3e1ad214898389ebc819, 256'h45da7b6fc8f4f766f82c5132735f2ed94130780b444e2e10c1484d5e45f64332},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{453, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h4589f0c24d1b2f89c2e806f667297c844c63330d6b9a079b2bdd2d95247e3eae, 256'h75daa1da09a3f1ed8de1aacc7039a721c46f9ebcd4672750f2fd9c2f70f1e6ed},  // lens: hash=512b(64B), x=232b(29B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{456, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h2f11d967790dd4387a218929b3fc0f130238ec6fd9321348fe631a1e607bd742, 256'h3b52a42606d0daa135092d89ab74b3c4e72b4ed213137406d4b50fa84c4ea049},  // lens: hash=512b(64B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{457, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h192d299e96272a0c49ed1b15f9047b54b4878eaf350a7b2f5439b1e3c83f9703, 256'h26513e9cbbaca7946f3d6d90b5cc65a985cdfe089734f944ab74842a4dc4127d},  // lens: hash=512b(64B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{459, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h37fd00b14ff469a8bb4d2f9c6ca228c4c24b85719389a46099653c41174e9afd, 256'h5f64dc68893cf3186df3e83af70e96e9f2103d25b8ddffecda96e8e9181619cf}  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
};
`endif // WYCHERPROOF_SECP256R1_SHA3512_SV
