`ifndef WYCHERPROOF_PACKAGE_SV
`define WYCHERPROOF_PACKAGE_SV
package wycherproof_pkg;

  `include "wycherproof_vectors/secp160k1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp160k1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp160r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp160r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp160r2_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp160r2_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp192k1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp192k1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp192r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp192r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha_224_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha_224_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha3_224_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha3_256_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha3_512_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp224r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp256k1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp256k1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp256k1_sha3_256_vectors.sv"
  `include "wycherproof_vectors/secp256k1_sha3_512_vectors.sv"
  `include "wycherproof_vectors/secp256k1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp256k1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp256r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp256r1_sha_256_vectors.sv"
  `include "wycherproof_vectors/secp256r1_sha3_256_vectors.sv"
  `include "wycherproof_vectors/secp256r1_sha3_512_vectors.sv"
  `include "wycherproof_vectors/secp256r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp256r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp384r1_sha_384_vectors.sv"
  `include "wycherproof_vectors/secp384r1_sha_384_vectors.sv"
  `include "wycherproof_vectors/secp384r1_sha3_384_vectors.sv"
  `include "wycherproof_vectors/secp384r1_sha3_512_vectors.sv"
  `include "wycherproof_vectors/secp384r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp384r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp521r1_sha3_512_vectors.sv"
  `include "wycherproof_vectors/secp521r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/secp521r1_sha_512_vectors.sv"
  `include "wycherproof_vectors/v1/secp256k1_sha_256_vectors.sv"

endpackage : wycherproof_pkg
`endif
