`ifndef WYCHERPROOF_SECP192K1_SHA256_SV
`define WYCHERPROOF_SECP192K1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp192k1_sha256;

localparam int TEST_VECTORS_SECP192K1_SHA256_NUM = 229;

ecdsa_vector_secp192k1_sha256 test_vectors_secp192k1_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 200'h009ecb5311ba692e0d41d5d7654d0c8c4ea7f71eb92b2e4996},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'hd781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{3, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{96, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 216'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a8140000, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=216b(27B), s=192b(24B)
  '{97, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 208'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f70000},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=208b(26B)
  '{101, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 216'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a8140500, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=216b(27B), s=192b(24B)
  '{102, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 208'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f70500},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=208b(26B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 0, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=0b(0B), s=192b(24B)
  '{118, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 0},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=0b(0B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h02d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6334acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a894, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b377},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a8, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 184'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=184b(23B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 184'h34acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=184b(23B)
  '{128, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 32976'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a8140000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=32976b(4122B), s=192b(24B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 208'hff00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=208b(26B), s=192b(24B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 200'hff6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=192b(24B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 32968'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f70000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=32968b(4121B)
  '{136, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h01d781b83e5846f00406b23fce604ca5b7606846f47c8fa5a1, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'hd781b83e5846f00406b23fd21266ad894195ba1f92d1aa87, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{138, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'hff287e47c1a7b90ffbf94dc02fc6a6565faf00ff75f84f57ec, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h287e47c1a7b90ffbf94dc02ded995276be6a45e06d2e5579, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{140, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'hfe287e47c1a7b90ffbf94dc0319fb35a489f97b90b83705a5f, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{141, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h01d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{142, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h287e47c1a7b90ffbf94dc02fc6a6565faf00ff75f84f57ec, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{143, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 200'h016134acee4596d1f2be2a289700d96bdf76db6e1bbe8fb184},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 200'hff6134acee4596d1f2be2a289ab2f373b15808e146d4d1b66a},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h9ecb5311ba692e0d41d5d76726199037988dd84eb64f4c09},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 200'hfe9ecb5311ba692e0d41d5d768ff269420892491e441704e7c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 200'h016134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 200'h009ecb5311ba692e0d41d5d76726199037988dd84eb64f4c09},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{153, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{159, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{163, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{169, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{176, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{179, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{180, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{182, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{183, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{184, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{189, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{190, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{192, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{193, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{194, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{195, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{196, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{199, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{200, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{201, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{202, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{203, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{204, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{205, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{206, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{209, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{210, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{211, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{212, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{213, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{214, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{215, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{216, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{219, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{220, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{221, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{222, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{223, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{224, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{225, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee37},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{226, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee38},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{238, 1'b1, 256'ha16c855ca4e25b5c5d4a588ef548fceb85f054765f64bfad874b67c415926488, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h0c9347bc9ee64533cd1a7825b5c4317f58b3c2d6d757ed8c, 192'h11ed5de0780eea59f2ad67a045e259f34208de10fd963ce5},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{239, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00db8557bc7915b9aec747bef876368ec13f8ba37f58a34c95, 200'h00823afc12256a13d24d6ec481eb673a5b5e58a4276e7dc401},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{240, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h4771aa9cd70dafe9c7dcccf139b5418bb626280a970b3163, 200'h00a23ea28ae4966a62d33f872b1379471828dd77ff89d211e8},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{241, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h008d60cad970bdaebf1e4031e7217c33840880310b2f4c3352, 200'h00977040c9b1b002b8f7474aac033a8aa3e5a665ac31e04c6e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{242, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00f15f1fd8acc9ff12877ea04f6caa8852445c80b3ec866124, 200'h00cd2ae16c50101eef38f878906acd2fd0a0a8e0622adb12c8},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{243, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h6ed69ce7626f0677cf82a1d4c9ffe1930cedcb6c0826c06f, 200'h00ec2347ff49bd92415f0731daaf73348631ce0dcb0b9d9034},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{244, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00a34cdbb418ad82a7a8e1fcf709e96bcc292d4c548995d3c1, 200'h00adcedd7ca763df0154f128901d23cae7c34df711966cc0da},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{245, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h3a4bf99959dbc04bca3ae3c8495bab859075c5ed793b8e6a, 200'h00e64279e29b46e8ff981573e145fc698a93529035d4f9a7f8},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{246, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h0099d169f6353e07bdfd2411c19d11b32848d86ffc87f2336e, 192'h29b1e44d5a3ae433d645cd19c6a59a7dab3b03b66a8730be},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{247, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00991d09d32e0815faa81611771897cebb8472c12c18fcc8e4, 200'h0091b6fa9d2cbf80b58304d4c3aafae5c200f3479c97e196bf},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{248, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h4b570cc266f484d1e18fbb4a4f9c9d67ded1c40fc1ae2e6a, 200'h00b3907e01b0c1b2248c025e3b7c70c9b43979d3148eb26190},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{249, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h25de156e669ab3310bcd79821ad5fb97333bfb26f5ba29a3, 192'h2deefd2ac3596fb1f17a3db7b17f2752daca453ea8fb177c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{250, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h4f9eb4f1b8be3bf608c91289d0ffa7281e2176bd04e2fb5c, 192'h694c480fb0b02edc9daa5006986ad96216fd673b277c8583},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{251, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00dbfef4abcdfc6c66cbe4c0940130fde5dc5323e80537a7e2, 200'h00c181d8297e962dcfd38c92c1687b54cb2d95002f05683a99},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{252, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00934db7759d0b26063f1b3fe9f69f4e2e363b700e67f6416c, 200'h00823dc4d2cb9473fed0cf7f884b48f067ec4686362840c442},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{253, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00b11eadceefb34b60728cafd6fc8aad2a6579df4a52b691f5, 200'h0083d6288af6908a1a861ac91b1eb84d8f26d878f73ef34159},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{254, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h1e1d9d3f3ff732612378e0fb564f5d80cabe7e4b7d37c464, 200'h00be5cf54130240da503be67579637e7f245efeb40523b48bd},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{255, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00fc1274b8e27dc06adb7ac57c06ab4d3aeca8632b611406b5, 192'h7b55e6637df8356001ffbd5fb2e36fb737b3a1ddf1b35b89},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{256, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h02debe93920d079a0f9239eac03fa5eb20788cf915982909, 192'h371d0950c7d32aef6e05ae5ce3e043cf9a129191897a60ab},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{257, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00f7936ca4c577a4e8fe1fdc406381b32f82cc4a523b7023b1, 192'h296f693ec6360effc49c43959bde6265625ab4bfc225ce79},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{258, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00e6a29c8032e75c5818f22760b4711cf0a5f8ea3aea1f3073, 192'h7285528eb3041ae6f630778e22ce4ae884fb0a38dc950ac5},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{259, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h008cb6072c12069e5b0e568855fc209a3cac9885228e464e0f, 192'h089932adcae5e75eac203c12c6e86f424fbf55a717d5ba72},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{260, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h01409e9e5dd41cf9e5eed02cca49c3584f7e26ee4508d244, 200'h00bb8af45b63c1a344c839f4ebc2e5fd6bcd484b7af15f4a47},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{261, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00f14781881a2687c3bcafb210c49572b80248f5f36492d3b4, 192'h368d5952265d5517ade8d638eb312b03c925e4234a27bda1},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{262, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h009ac57b79055eee9ced09ac450aa0b84efe94fef74a40d9bf, 200'h00da4f41332b79a46ffb811ff10ca443ff5cee330143c2c6d0},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{263, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h727c6a44c692934be6e761f1bf89b436ec37c5e80c7560c1, 200'h009eedd523f8e01e635743a2b64619ac4c3e34d63831dda18b},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{264, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h48ad2b9451c5a6bffaff95874dd0e8000870df00c89ef274, 200'h00d7d59fea2ad4c5688c26037f89f0b8d883eb546f58433cc7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{265, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h2b6a95e8a60194d2d850f510b35120c7eb454a52dc2f92f9, 200'h00ffb706d807e6e4bcfd89e9b696ebe233c62c10a301c54858},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{266, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h2a70e9a299ecc9cd6490ecf263018b1aef248fef4bdb92b3, 200'h00c1599dac7241f8d1c630cda9a53eef1e87cf5b7178845f0a},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{267, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h36960dea8d79e3239d9c84d26f45982726801d7367f4aff8, 200'h00be23a608dcefe3c7409978b2cb8549227e2286ecb538c0ca},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{268, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h1da1bd31f9aebdb4da362f892ce9594450ba808e8ed5a561, 192'h46d7556ce3d34ef78c0a6ec454c4cae1d4464247bfe007c5},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{269, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h54bbc9994c16eaec46aaca95a703d374e91025bd6bac5676, 192'h6671ff343c58fa6a965cb0ed66090a0e3ff2ee9287dc6d13},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{270, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00a778cac2653046d0bef2cadb79cf24d588154ff35fb771d8, 192'h6a534b96ea6e4dbe1216db94a6132767d529102d94e7a944},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{271, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00992969b923959673afa12cad8578fb8067b6771b3f7fc2d8, 200'h00d1c3dedc0ce64f83f5ef56a5be20bddb2429902f929e245b},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{272, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00caabe0ebec465309b3a7802f8e95a209650f32ff74d6656a, 192'h34e40a8b6caaa063b03f72b000deaaeca5002e3d3efd6065},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{273, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h05f6b01f861391aa3326218df2cf89c572e65ef7beb4d241, 200'h00c9792f3cbe70ebd5e8a3566ae8344a58484305152eb6cfcc},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{274, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h0438234511040ff052fa84f15a43022f926bb706821d3be3, 192'h7e85ed42bca80d528c1b6b981677fd2ab353a81a096fbb87},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{275, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h448683d5003b466baf2c373da244a58125bb649afe14fae3, 200'h00ba251ba99f8f8624580aa19e5585cac19bc9eff5fc078367},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{276, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h009c827ab885ab43e809db2dd881a1141e0d13762c67167c25, 200'h00e60f0185e26ef8c5030eb1f9173beb9f38e4d35157239394},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{277, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h4ae9a2f972b71b2883862d69db9061bd1f7c47ae003e46a7, 192'h31ee553e8940621d8724103e3ce080dfab61b0c51f466da4},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{278, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h0080acd9c4aed0f5b5884cf50c0f2bb322c9445c0ed8e4cd12, 192'h08cddedf81c5c5fba6c42ccddd1f55a907a63621469e2822},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{279, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00f724abbec061bc29b6b2d3a370281e4d56b0225244ceb8fb, 200'h00c80009ce8d87d8988c305d8a69bbf37a7d3f0b1e72f3444b},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{280, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h0094d3d2ac3e34ba421fe919e3326837a29efeae4660809806, 192'h71c1a1dff0dc627b18c39e50634e0bd31969163e976cdf76},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{281, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h50892f46b087ce202c39cbade6f3ac5d344d3a9b1cbae513, 192'h37bc179d7aa0cdd36c479df175d8968630e0875cb84567d6},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{282, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h6ca8a34e1ad10e46abf3ef5a7d8b94c0de703611c4e8e0e8, 200'h00adc1a44bed4bf73a47b11fa72689ba9f63275be4911ba360},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{283, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h1fde9536082e359e2e930e2d43e364cc62493385623510cc, 200'h00bd5c6e0f8f573e60f3ca1b7ab29a112c50e355bc9beb02ee},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{284, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00ad83df6dec32487c9ccebec2f98f335c4e889bcf573db16c, 192'h7d84f6b32a7ea7e78eef051e626cb34b183d96c16d918b00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{285, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h67534cebf5736c79df01a83d6d67d6e757f496cc14ecb60d, 200'h00c84db7860a115eb0215a412fab9575ca9971fe4e3a13c0bc},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{286, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00850f2891e3b3874a2de647ce777504069eae5af18e64d3ce, 200'h00c7f0973f4433bbcb1974250af73cb124d2e559afa91101ba},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{287, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h008e1c922ef2d3d16ac6830e0db5f16f6ca9fd680991600a92, 192'h644d5c24b90a9dcbf2fa9cd15a2aab2f0a189b97a7360477},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{288, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00ce211ee377411353e62b7d07159ba7080a890accf9b185d1, 200'h00ee03f5d17b54ce1ba4d7e44a4b5344a44ee3588988a9909d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{289, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00e591fb2afdd2250a6543ae797ba7b4b863b0b1186afb2ec4, 192'h1f59d7c39b4cb9281602fee77d677743f26ec6842e4e7b53},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{290, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h1838557c794373b31602d065a36853486b2c501d53004294, 192'h388eb4817ef3b2273563cb07afdce8ae19c6aa9b78d8d7ac},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{291, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00b55b6effb9a94eb81dc11cb1efb213dee62bf466d165b75a, 192'h4b6b456f24387db822d9c9b7965e3d835237ea78565ce95f},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{292, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h57f4795eda4e8ce0cc7447f65b1c63938c171126dceb3fe3, 192'h277c0487e82b8f3bbc8d320be12a5ee8ebf29544577cd146},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{293, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 200'h00c53070be8227256e660d9ca572062d2dde4be55befefe58d, 200'h00c30fc40af6fa6f84f3219e72a52ec295b7f94417e67c6e6d},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{294, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h70779f44a7711a14cc2a732870c969c9fc3eae11727727a7, 200'h00f83f576bd9347b4918bd5333eb4d93a285e71f4fa86dc409, 104'h01d90d03e8f096b9948b20f0a9, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8a},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=104b(13B), s=200b(25B)
  '{295, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h70779f44a7711a14cc2a732870c969c9fc3eae11727727a7, 200'h00f83f576bd9347b4918bd5333eb4d93a285e71f4fa86dc409, 200'h00fffffffffffffffffffffffffffffffffffffffeffffee36, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8a},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{296, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h1937a518d51769dd68a57973b2fb4cf342eea3449458646c, 192'h2e688800bca2ba941874b5a88ff09b757a408a5b09d8474b, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8b, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8a},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h008be871c72c4a0b3fc37d0a50401fd3b968dc2eab13bd3696, 200'h00d4e571d5bb93193ade7cfb88cfc50974227b8473f008dc41, 192'h7fffffffffffffffffffffffffffffffffffffffffffffff, 200'h00da23d70c4ab11a41d6b4578b5360b607ab913b00c36b4520},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5d9a58ab6292a92b6d7e050f90094e09a3bb38f98fb331aa, 200'h0084c8afb5a6a68fae7e23971efccd15e631c8405509814fa5, 192'h7fffffffffffffffffffffffffffffffffffffffffffffff, 200'h00d767f661ddab5ab0432826fa4da22e596839f8f25fb2d50d},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h6e7ada341f8d180bca044695af5394e3380164233cf9764e, 192'h00a893be62c1b460767f412761d2053bd49eaf549df1cf47, 8'h01, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7c0c136b0b58d9c1b8adaa1a2d7b4bbfa67f485ba258e6dc, 192'h56f829f77d6bee7f02bb0b1b0b628337be66d83656eac152, 8'h01, 8'h02},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4a352661886a1ff22d1376abf349caea36ada82e7856c77b, 192'h6bafd111064272ade6c396c584f857b4801a5547702f4278, 8'h01, 8'h03},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{302, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4a352661886a1ff22d1376abf349caea36ada82e7856c77b, 192'h6bafd111064272ade6c396c584f857b4801a5547702f4278, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd8e, 8'h03},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0f73a6dd1b1193defca5b3372c783c7938553e8f8251eab0, 192'h5985e813887dca413b082db9ed640854d916f1fd598ffff8, 8'h01, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74f1d414},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=200b(25B)
  '{304, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0ac0601e26e29f23f6de5a71e6ac2473d7d5c8018c04a2b5, 200'h00f0987bf80c7954f9211c3acf7ca23a0039800c523ac2970f, 16'h0102, 192'h1a3468d1a3468d1a3468d1a31620ef794a24fb1d09f28ad6},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=16b(2B), s=192b(24B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h1c0c3e57759ffe70a11d5be9955cc5593882fe7cae23b168, 200'h00c1bc39cdc60d3156c04acc5b8565ed8407c251e9e1ff3485, 56'h2d9b4d347952cc, 200'h00ae8a60731be897b57fae4ace724ea52f89cc05ae6a3e68e3},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=56b(7B), s=200b(25B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h53c62f3128456bd96b1c7b95c591ff4cda4332b0d54d0629, 200'h00e561307a73f26f12179b9cfd6304c07c6ec261b8d08243a9, 104'h1033e67e37b32b445580bf4efc, 192'h28d728d728d728d728d728d6dd5f8ad4dc9b410606b10596},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=104b(13B), s=192b(24B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h61e6de690644cc59228a7fb723f4233b3615b7285c3caef3, 192'h113ea0243966be0e19f146b24efe7d812e7c80033fa8a03d, 16'h0102, 192'h18e328c9b6a27246966d675cccdb4c300f4b029466ee5b79},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=16b(2B), s=192b(24B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h008637d3b364384b999e82460b12660029fb8d72e2e47b9eae, 192'h41d8e59ab0ac5df6feb34639438b1ed4da2a7c3ebcd72cf8, 104'h062522bbd3ecbe7c39e93e7c25, 192'h18e328c9b6a27246966d675cccdb4c300f4b029466ee5b79},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=104b(13B), s=192b(24B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h572974ebd982bc0a38f6546a347745b7a071c4d6333fee43, 200'h00a78c487f6ffc4810d480c9c6086a0c9f8f2385e77cd9279e, 200'h00fffffffffffffffffffffffe26f2fc170f69466a74defd0e, 192'h555555555555555555555554b7a65407afcdc2237c4a5484},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0a03d1b9b71bfb929ccc2f93f0f22ccd012679ac7517509d, 192'h3425a86e0982e15e4a012d9810693a6ca1647175f1d3a125, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=8b(1B)
  '{311, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0a03d1b9b71bfb929ccc2f93f0f22ccd012679ac7517509d, 192'h3425a86e0982e15e4a012d9810693a6ca1647175f1d3a125, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h3ebe178e893f584ff15c5eaf86fae4221f1de334834b6625, 192'h318e73821c2d63c0289171e0a0bc702542ed4ae0c6662395, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec6, 192'h555555555555555555555554b7a65407afcdc2237c4a5484},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{313, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h008e6a351293a941095f3ead178835f38507a108c5facfdf84, 200'h00b16293ba6f5d5ad63e3bb977ee7ad50cdbbb6a8f4602aac2, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec7, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec6},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h008030f67279e1099e19b1a54ebe8e6945620b10b476925d14, 192'h2a28bda0e6cb2bd718e9e87fb2b5441c38347a2c3a0146ed, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec7, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec7},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{315, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0091185b730be9b119fad97d216164b3af07fbb217d4c337ce, 192'h436fd95c99b7f0df881b0586c707b4c67fb89e373a219ad2, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 200'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c88},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h321a763b434b23fee5ee41b369fd48f4a5b64df73fcad9ea, 200'h009340d92cd1f67d75393be503fcace7212876b71f4c717996, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 192'h44a5ad0bd0636d9e12bc9e0892d05a340f325ea749b7f105},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c579dce46d22d891fa2fd06e3f8e2d0664f5f040ae42a78c, 192'h483e6407c797bfe22dcb09a66a5564b6a82120c130a130e0, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 192'h555555555555555555555554b7a65407afcdc2237c4a5484},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5b6ed27bc9e836b8027a62e1e6d42c8478b6532e93fdb12a, 200'h00f7d82a16221b613662c8b62d6507fa1185526174209f15dd, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 200'h00aaaaaaaaaaaaaaaaaaaaaaa96f4ca80f5f9b8446f894a909},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00898b80717733e395dfdca2d7135fce6a9cb422ea902314a7, 192'h4420d6419551c2d5a49898a02ab409cb855a62bf4853de08, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h0093c8c651653430cb4f1675fbe90734a8afe00f648aacae07},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d51b0f873aab3e12fcf2595df0ca3b0184e2035d5b3b3e72, 200'h00d49ccc303545f1d6747faa50d6258d55336c85f31e9db2e0, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h5609ac29f2adf8f19445587a7b083b200127623c11a53fb7},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e461f50514aa00e42cf2a3843c95c5e6198fb62c16da2be7, 192'h46e935ed8899edf7fb8c7f880a439b89c9721293bc3a1ec5, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h0097614ee6f88e6a88648d43ab92c20bdc3f074eacbb26d47d},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e3c17e3321bbf47cd866a640e56d9f30440a1170b0b35dea, 200'h00945c871de164867b50b8f44153c35d549a09210d3efc7096, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h0dcf2f2634c548a744a5ad0bb6deebc51800e1ecf4ab5a57},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h506735ecbb1df64bc52226815a323195f79c2d4e7d398c76, 192'h0c81460c20101ffc243a42a2c618088896c7826b7c8d40d8, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00f2f2634c548a744a5ad0bd0475ebadaecfa64bce46038ad4},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00854119117aa43693035af1736f8095e3d3fac40d39a3d5db, 200'h00e83f70ccb798e9b9db84a959dddf6b99c575dd9576ead5a7, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00e5e4c698a914e894b5a17a0ac4e45f468fe351321728181b},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00acc7b989fcf4270cf688bb12e1a9a98e320a194ae0a9f938, 200'h008537068f16aa3c575f189df9be197a7dec4ff7f2f736cf9b, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h34c548a744a5ad0bd0636d9db1396bf8ff1987e588567a12},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4112a1eb92dc6f34e4ce23290b9469728f1c74f495a2b664, 200'h00900900d77fa23e99dca9e3015e5b34cd5e5035cb86bc3730, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00a8d472a340c9c2545f8e65efcfbabf922ae645c50ebef1b2},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{327, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h3a107a26b2798afc115ca9cf473b801ab5388415cdd07d42, 192'h7c815c7b542d09d621be6c9e6ef299c4e1d65748b0665400, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h008f47ba72d653756936634785f0f78dafcc48fa3f3bca2d69},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4f911c19941d1628a75335d80e34dcd59c59b46ec0e7a703, 200'h00a70701af5a67581953b5b406b65c245e6f1137ab63199a66, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h361b9cd74d65e79a5874c5011ef5e3b72fc49b82f51927c3},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009504d8916295ee0e37028cf98b4ac4695fc5d9169c22c39f, 200'h00d1dd393e76f50871c9a8ec3d381cbcef14d1ae57396a7aff, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h6c3739ae9acbcf34b0e98a023debc76e5f893705ea324f86},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00a75790f8ef02dc29cfb095fffe450e9de57a85c3e09b0e20, 200'h00bf02919d1af324098da7731a3bacc5bb71eee7ab24ad8ff4, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00a252d685e831b6cf095e4f035ce1ab258f4dd288df4b7749},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h565b7b8da8bd1dfde987d73b3037b6b0c22f0f03ba526f38, 200'h00ea50fa9fbf19711b04a46b9fe30032f4215cc72b70f32b4e, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00cbb0a7737c4735443246a1d4dcda83f9a7384a8b9802e905},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{332, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00da8fa3039de9c6d080640cc63bb80546f2c60bc4109ee3fd, 200'h00ff6b94e7f86cc4b9d9c5202823af1c989d6f34686d1d85c4, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00d5555555555555555555555419f752ba0a462ef1a33f53b2},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h00e3ebcc961c21e5377993a6ae56169cfb02b6b29fada4fe, 192'h12a947f948c11cb04f5349e7eab3de4db904359ea41e7b11, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h71947adb1fecb13a7be2f9587ab6d22e2b88223d145b2948},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{334, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h025c53fea2b2e10175f2887693241e7271b308510a479721, 192'h750ba51102b54f2a4bb10f6033c8792415665b85f88c88dc, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00e5f84a7d49e369ab1469d151beec3e137ffbce835a1e3d76},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{335, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00b645468ca1107a766387231b4be740698b3468f1de6ca6e7, 200'h00d3a83176c30b7cccf7feb6c1e299c28b1f2fcb891125abe7, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h080f8ea15811caeb7ffffffff11ad88e21bd2c3dd7e6f462},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h572b205771aa8a4bd40980103ce547e11066b75c9c98a926, 200'h00be118a6763d86738075ee9c757b1756c7acd453ad6d5db4f, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00f8ea15811caeb7fffffffffe340ad6941e20a843ffc75980},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{337, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009e8fb05735832aa74f3546ca43fb91dd6876c2fa773851d7, 192'h2dee0143e2446bf9bbd7779f6fce9d6ae0938832dca2cba6, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00f1d42b02395d6ffffffffffe4122b1112cd80a1d8aafb573},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7e1e836b005fec913626163c76a4be541a2461842975ab36, 200'h009b08b9786438ddfc226586479ad7f6b1bc4a8ce57b33e8fb, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h5811caeb7fffffffffffffff5d42a5d24dbecd9d8bdb5453},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{339, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h109224c4593360afcc68b9657351c2547ebf8e6eb9529171, 192'h5901934cde484511c3a0927888fab4279898b5b1d2fd2418, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h35f5f5f5f5f5f5f5f5f5f5f58fee224b3f8f2d4e2d4931ab},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{340, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5311d7f38eedd5802452075949558664fc85dd38917490fe, 192'h6a7e77e633b1886ca2df3b0b96e9cf9d935710fd71d19f7d, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00e1af286bca1af286bca1af26c48890b651284c7a32ac9205},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h46104a66f225bc3bfba7e6e55774dbaa7b8d4f35bd046dfe, 200'h00dafd7c2a12a3ca7d84229073a6dffc5dd2fe961e00836e7f, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h0095555555555555555555555419f752ba0a462ef1a33f53b4},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{342, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009816a33b6358273f3a9ecb25c0587c7f75cc6b6261a62f19, 192'h3a0d01b21b285109264df65d0ab2f4dc9e8a728e02955c44, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h2aaaaaaaaaaaaaaaaaaaaaaa0cfba95d05231778d19fa9db},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{343, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cac32981b0eebd5641bb9118d6f3ab2ecbc1ec90182e0798, 192'h363a02c11e577a366058830ff90f88a1fe2f2e380e23adbf, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 200'h00bffffffffffffffffffffffe26f2fc170f69466a74defd8f},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{344, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7ed480fc2ae377d350f1e89cc704810522bd1010529debe7, 192'h343c9ae0ee77f6737c874565346417d26d99e295474d46af, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h72fc253ea4f1b4d58a34e8a8df761f09bffde741ad0f1ebb},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{345, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00a92126a3121c77cc9d36c071e5d25dd777cb0751eea960d0, 192'h332ab2bde6590c6e0fd6c2068d384da997e6274fbfd5bd06, 192'h4ca731ee2d7eac575784526b77c25003b24e72d5084d8456, 200'h00a12629aae1c4360c7e560c0c0188d09171bfb620215e08a0},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{346, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00a92126a3121c77cc9d36c071e5d25dd777cb0751eea960d0, 200'h00ccd54d4219a6f391f0293df972c7b2566819d8af402a3131, 192'h4ca731ee2d7eac575784526b77c25003b24e72d5084d8456, 200'h00a12629aae1c4360c7e560c0c0188d09171bfb620215e08a0},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{347, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00fb2b20bfa7a9925006623c5380d6870a9ffc1151eb54919c, 200'h0081bc177fe523ce4a89170e8b03680132d6911dc6d154c329, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 192'h333333333333333333333332d496ff37cfe1dae2175fcc4f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{348, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h46214be9f3858d360a22f8e5d367c2461b542167364aed54, 200'h00ba162fdf946fa2da9175b61c98ed89402d8ce3744e0175b0, 200'h00f091cf6331b1747684f5d2549cd1d4b3a8bed93b94f93cb6, 192'h555555555555555555555554b7a65407afcdc2237c4a5484},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d9c3df86bcd75a2134357cd6171732414be030f454b87266, 200'h00efb71c8bdb526a9238fabaefbfdc240ba86a1f315cb99773, 200'h00f091cf6331b1747684f5d2549cd1d4b3a8bed93b94f93cb6, 200'h00b6db6db6db6db6db6db6db6c64f6b41078b8e927780cfe40},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7aa940cae4ac1f9f3b2ca8826541c5d9028c3374199c0b38, 200'h00d38821fa104f582a779cc4eecfba28984df1cd52c1bf7133, 200'h00f091cf6331b1747684f5d2549cd1d4b3a8bed93b94f93cb6, 200'h009999999999999999999999987dc4fda76fa590a6461f64ee},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h74393ae3827d99146c93121e09f20c8abeef24a0df3aa24d, 200'h008a0c78af68f0cbce09ceb71011be5b1a67b653b5ca5a9e65, 200'h00f091cf6331b1747684f5d2549cd1d4b3a8bed93b94f93cb6, 192'h666666666666666666666665a92dfe6f9fc3b5c42ebf989f},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0082236bca1130e814226ebdc51ceef77b12f0acf75529209c, 200'h00d2b2e825b5eed059a8b284c768b2ca887951a6bacec7b505, 200'h00f091cf6331b1747684f5d2549cd1d4b3a8bed93b94f93cb6, 192'h492492492492492492492491c1fc480696b05d42fcd1ff4d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5eb0103ffd191c7e743328eadf65d5e0d111f49cf7d5fb8b, 200'h00dda35a625496a8007877a0b40632930402bdb09767cd218d, 200'h00f091cf6331b1747684f5d2549cd1d4b3a8bed93b94f93cb6, 192'h0eb10e5bb837a2b8056c361dad570a9ed7e4d14114fe6e0e},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h1b29886ffb76447b05b19dc3b30d38dee455135026da8357, 200'h00bde5d4d6400488c764411ec39e78a58a1d22789e33459114, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 192'h555555555555555555555554b7a65407afcdc2237c4a5484},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ce38eb489f4791ba70216d25a97039fa1c29ef0347fcc85a, 200'h00dbf1a45428550a6de645b0796d4ec33e73174998b1dd3944, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 200'h00b6db6db6db6db6db6db6db6c64f6b41078b8e927780cfe40},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ec2b5ce564ddb6785c7687d1e1297a066b8cef67911e31f2, 192'h6e0f2c5ad2cf95b2753d7de9ebb5ff0d6bb95455de865488, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 200'h009999999999999999999999987dc4fda76fa590a6461f64ee},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00acbeb945f5a6ec5a6f944df4688a6d38f2995db3089918eb, 200'h00f2b5e522a97baf3e6afacbca779ebe06665e6390bb88f950, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 192'h666666666666666666666665a92dfe6f9fc3b5c42ebf989f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00b7c68007cc4017c7787c4beec984252eebaf57f4b699f003, 200'h00c1d8daa7a0312ec4de5afa5024f5762fa2da773800963018, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 192'h492492492492492492492491c1fc480696b05d42fcd1ff4d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7d7c2fa76599eaf664ddd75c7ab1ea7deb5191eb3327c48b, 192'h78c029886e4467b49adc5460fb7ad6facf5a2902bb1c0974, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 192'h0eb10e5bb837a2b8056c361dad570a9ed7e4d14114fe6e0e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{360, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 200'h009b2f2f6d9c5628a7844163d015be86344082aa88d95e2f9d, 200'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c88, 192'h249249249249249249249248e0fe24034b582ea17e68ffa6},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{361, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 200'h009b2f2f6d9c5628a7844163d015be86344082aa88d95e2f9d, 192'h44a5ad0bd0636d9e12bc9e0892d05a340f325ea749b7f105, 192'h249249249249249249249248e0fe24034b582ea17e68ffa6},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{362, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 192'h64d0d09263a9d7587bbe9c2fea4179cbbf7d557626a1be9a, 200'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c88, 192'h249249249249249249249248e0fe24034b582ea17e68ffa6},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{363, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 192'h64d0d09263a9d7587bbe9c2fea4179cbbf7d557626a1be9a, 192'h44a5ad0bd0636d9e12bc9e0892d05a340f325ea749b7f105, 192'h249249249249249249249248e0fe24034b582ea17e68ffa6},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{364, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 192'h04a4e7bedc7d8137aade86c1a4d223ad704e63dad4717c49, 192'h3efc196def1cad9823c91f6b8be2611164b93cca4bb2c559, 192'h5ca564801c724e9027e6d39f006ec3f63bd8d3829fdd7850, 192'h6eaec4b21473db322e9924f12d2a260467c0ed58882e7134},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{365, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 192'h04a4e7bedc7d8137aade86c1a4d223ad704e63dad4717c49, 192'h3efc196def1cad9823c91f6b8be2611164b93cca4bb2c559, 192'h546e7cfe5f660f10a02cefdcb4bb4e0cc7a9fd43cc9e443f, 200'h0086d3a935dd62d5db7101e128f3f6048c490072a49a5ef047},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{366, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h04a4e7bedc7d8137aade86c1a4d223ad704e63dad4717c49, 192'h3efc196def1cad9823c91f6b8be2611164b93cca4bb2c559, 192'h4e64634ce6163b98ab39d573698ea05620721f389fc27da7, 200'h00df079942bb819f533a629945c970134d1017e8ae8ede25da},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{367, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 192'h04a4e7bedc7d8137aade86c1a4d223ad704e63dad4717c49, 192'h3efc196def1cad9823c91f6b8be2611164b93cca4bb2c559, 192'h28d91785c005c416c436222a06578939d12c9ead1cfcd63c, 200'h00828921b3e632424caa08ce947d2ef43a3b9ccb89f5a74820}  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
};
`endif // WYCHERPROOF_SECP192K1_SHA256_SV
