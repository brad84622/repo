`ifndef WYCHERPROOF_SECP192K1_SHA256_SV
`define WYCHERPROOF_SECP192K1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp192k1_sha256;

localparam int TEST_VECTORS_SECP192K1_SHA256_NUM = 56;

ecdsa_vector_secp192k1_sha256 test_vectors_secp192k1_sha256 [] = '{
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'hd781b83e5846f00406b23fd03959a9a050ff008a07b0a814, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 0, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=0b(0B), s=192b(24B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h00d781b83e5846f00406b23fd03959a9a050ff008a07b0a8, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=192b(24B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'hd781b83e5846f00406b23fd21266ad894195ba1f92d1aa87, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h287e47c1a7b90ffbf94dc02ded995276be6a45e06d2e5579, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{142, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h287e47c1a7b90ffbf94dc02fc6a6565faf00ff75f84f57ec, 192'h6134acee4596d1f2be2a2898d9e66fc8677227b149b0b3f7},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h00, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{159, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'h01, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{169, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 8'hff, 8'hff},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{238, 1'b1, 256'ha16c855ca4e25b5c5d4a588ef548fceb85f054765f64bfad874b67c415926488, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h0c9347bc9ee64533cd1a7825b5c4317f58b3c2d6d757ed8c, 192'h11ed5de0780eea59f2ad67a045e259f34208de10fd963ce5},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{249, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h25de156e669ab3310bcd79821ad5fb97333bfb26f5ba29a3, 192'h2deefd2ac3596fb1f17a3db7b17f2752daca453ea8fb177c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{250, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h4f9eb4f1b8be3bf608c91289d0ffa7281e2176bd04e2fb5c, 192'h694c480fb0b02edc9daa5006986ad96216fd673b277c8583},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{256, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h02debe93920d079a0f9239eac03fa5eb20788cf915982909, 192'h371d0950c7d32aef6e05ae5ce3e043cf9a129191897a60ab},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{268, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h1da1bd31f9aebdb4da362f892ce9594450ba808e8ed5a561, 192'h46d7556ce3d34ef78c0a6ec454c4cae1d4464247bfe007c5},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{269, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h54bbc9994c16eaec46aaca95a703d374e91025bd6bac5676, 192'h6671ff343c58fa6a965cb0ed66090a0e3ff2ee9287dc6d13},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{274, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h0438234511040ff052fa84f15a43022f926bb706821d3be3, 192'h7e85ed42bca80d528c1b6b981677fd2ab353a81a096fbb87},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{277, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h4ae9a2f972b71b2883862d69db9061bd1f7c47ae003e46a7, 192'h31ee553e8940621d8724103e3ce080dfab61b0c51f466da4},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{281, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h50892f46b087ce202c39cbade6f3ac5d344d3a9b1cbae513, 192'h37bc179d7aa0cdd36c479df175d8968630e0875cb84567d6},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{290, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h1838557c794373b31602d065a36853486b2c501d53004294, 192'h388eb4817ef3b2273563cb07afdce8ae19c6aa9b78d8d7ac},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{292, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 192'h657a69e8020565f6bb0a6254d24e06805c75b6f1ad819d8c, 192'h490866832f75cb6fbb7427eee4d89a767fdd5065000300f9, 192'h57f4795eda4e8ce0cc7447f65b1c63938c171126dceb3fe3, 192'h277c0487e82b8f3bbc8d320be12a5ee8ebf29544577cd146},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h6e7ada341f8d180bca044695af5394e3380164233cf9764e, 192'h00a893be62c1b460767f412761d2053bd49eaf549df1cf47, 8'h01, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7c0c136b0b58d9c1b8adaa1a2d7b4bbfa67f485ba258e6dc, 192'h56f829f77d6bee7f02bb0b1b0b628337be66d83656eac152, 8'h01, 8'h02},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4a352661886a1ff22d1376abf349caea36ada82e7856c77b, 192'h6bafd111064272ade6c396c584f857b4801a5547702f4278, 8'h01, 8'h03},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{304, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0ac0601e26e29f23f6de5a71e6ac2473d7d5c8018c04a2b5, 200'h00f0987bf80c7954f9211c3acf7ca23a0039800c523ac2970f, 16'h0102, 192'h1a3468d1a3468d1a3468d1a31620ef794a24fb1d09f28ad6},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=16b(2B), s=192b(24B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h53c62f3128456bd96b1c7b95c591ff4cda4332b0d54d0629, 200'h00e561307a73f26f12179b9cfd6304c07c6ec261b8d08243a9, 104'h1033e67e37b32b445580bf4efc, 192'h28d728d728d728d728d728d6dd5f8ad4dc9b410606b10596},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=104b(13B), s=192b(24B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h61e6de690644cc59228a7fb723f4233b3615b7285c3caef3, 192'h113ea0243966be0e19f146b24efe7d812e7c80033fa8a03d, 16'h0102, 192'h18e328c9b6a27246966d675cccdb4c300f4b029466ee5b79},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=16b(2B), s=192b(24B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h008637d3b364384b999e82460b12660029fb8d72e2e47b9eae, 192'h41d8e59ab0ac5df6feb34639438b1ed4da2a7c3ebcd72cf8, 104'h062522bbd3ecbe7c39e93e7c25, 192'h18e328c9b6a27246966d675cccdb4c300f4b029466ee5b79},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=104b(13B), s=192b(24B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0a03d1b9b71bfb929ccc2f93f0f22ccd012679ac7517509d, 192'h3425a86e0982e15e4a012d9810693a6ca1647175f1d3a125, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 8'h01},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=8b(1B)
  '{311, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0a03d1b9b71bfb929ccc2f93f0f22ccd012679ac7517509d, 192'h3425a86e0982e15e4a012d9810693a6ca1647175f1d3a125, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 8'h00},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h3ebe178e893f584ff15c5eaf86fae4221f1de334834b6625, 192'h318e73821c2d63c0289171e0a0bc702542ed4ae0c6662395, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec6, 192'h555555555555555555555554b7a65407afcdc2237c4a5484},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{313, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h008e6a351293a941095f3ead178835f38507a108c5facfdf84, 200'h00b16293ba6f5d5ad63e3bb977ee7ad50cdbbb6a8f4602aac2, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec7, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec6},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h008030f67279e1099e19b1a54ebe8e6945620b10b476925d14, 192'h2a28bda0e6cb2bd718e9e87fb2b5441c38347a2c3a0146ed, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec7, 192'h7fffffffffffffffffffffff13797e0b87b4a3353a6f7ec7},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h321a763b434b23fee5ee41b369fd48f4a5b64df73fcad9ea, 200'h009340d92cd1f67d75393be503fcace7212876b71f4c717996, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 192'h44a5ad0bd0636d9e12bc9e0892d05a340f325ea749b7f105},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c579dce46d22d891fa2fd06e3f8e2d0664f5f040ae42a78c, 192'h483e6407c797bfe22dcb09a66a5564b6a82120c130a130e0, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 192'h555555555555555555555554b7a65407afcdc2237c4a5484},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d51b0f873aab3e12fcf2595df0ca3b0184e2035d5b3b3e72, 200'h00d49ccc303545f1d6747faa50d6258d55336c85f31e9db2e0, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h5609ac29f2adf8f19445587a7b083b200127623c11a53fb7},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e3c17e3321bbf47cd866a640e56d9f30440a1170b0b35dea, 200'h00945c871de164867b50b8f44153c35d549a09210d3efc7096, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h0dcf2f2634c548a744a5ad0bb6deebc51800e1ecf4ab5a57},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00acc7b989fcf4270cf688bb12e1a9a98e320a194ae0a9f938, 200'h008537068f16aa3c575f189df9be197a7dec4ff7f2f736cf9b, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h34c548a744a5ad0bd0636d9db1396bf8ff1987e588567a12},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4f911c19941d1628a75335d80e34dcd59c59b46ec0e7a703, 200'h00a70701af5a67581953b5b406b65c245e6f1137ab63199a66, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h361b9cd74d65e79a5874c5011ef5e3b72fc49b82f51927c3},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009504d8916295ee0e37028cf98b4ac4695fc5d9169c22c39f, 200'h00d1dd393e76f50871c9a8ec3d381cbcef14d1ae57396a7aff, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h6c3739ae9acbcf34b0e98a023debc76e5f893705ea324f86},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h00e3ebcc961c21e5377993a6ae56169cfb02b6b29fada4fe, 192'h12a947f948c11cb04f5349e7eab3de4db904359ea41e7b11, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h71947adb1fecb13a7be2f9587ab6d22e2b88223d145b2948},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{335, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00b645468ca1107a766387231b4be740698b3468f1de6ca6e7, 200'h00d3a83176c30b7cccf7feb6c1e299c28b1f2fcb891125abe7, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h080f8ea15811caeb7ffffffff11ad88e21bd2c3dd7e6f462},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7e1e836b005fec913626163c76a4be541a2461842975ab36, 200'h009b08b9786438ddfc226586479ad7f6b1bc4a8ce57b33e8fb, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h5811caeb7fffffffffffffff5d42a5d24dbecd9d8bdb5453},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{339, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h109224c4593360afcc68b9657351c2547ebf8e6eb9529171, 192'h5901934cde484511c3a0927888fab4279898b5b1d2fd2418, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h35f5f5f5f5f5f5f5f5f5f5f58fee224b3f8f2d4e2d4931ab},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{342, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009816a33b6358273f3a9ecb25c0587c7f75cc6b6261a62f19, 192'h3a0d01b21b285109264df65d0ab2f4dc9e8a728e02955c44, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h2aaaaaaaaaaaaaaaaaaaaaaa0cfba95d05231778d19fa9db},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{344, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7ed480fc2ae377d350f1e89cc704810522bd1010529debe7, 192'h343c9ae0ee77f6737c874565346417d26d99e295474d46af, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffc, 192'h72fc253ea4f1b4d58a34e8a8df761f09bffde741ad0f1ebb},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{347, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00fb2b20bfa7a9925006623c5380d6870a9ffc1151eb54919c, 200'h0081bc177fe523ce4a89170e8b03680132d6911dc6d154c329, 192'h555555555555555555555554b7a65407afcdc2237c4a5484, 192'h333333333333333333333332d496ff37cfe1dae2175fcc4f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{361, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 200'h009b2f2f6d9c5628a7844163d015be86344082aa88d95e2f9d, 192'h44a5ad0bd0636d9e12bc9e0892d05a340f325ea749b7f105, 192'h249249249249249249249248e0fe24034b582ea17e68ffa6},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{363, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00db4ff10ec057e9ae26b07d0280b7f4341da5d1b1eae06c7d, 192'h64d0d09263a9d7587bbe9c2fea4179cbbf7d557626a1be9a, 192'h44a5ad0bd0636d9e12bc9e0892d05a340f325ea749b7f105, 192'h249249249249249249249248e0fe24034b582ea17e68ffa6},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{364, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 192'h04a4e7bedc7d8137aade86c1a4d223ad704e63dad4717c49, 192'h3efc196def1cad9823c91f6b8be2611164b93cca4bb2c559, 192'h5ca564801c724e9027e6d39f006ec3f63bd8d3829fdd7850, 192'h6eaec4b21473db322e9924f12d2a260467c0ed58882e7134}  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
};
`endif // WYCHERPROOF_SECP192K1_SHA256_SV
