`ifndef WYCHERPROOF_SECP256R1_SHA3256_SV
`define WYCHERPROOF_SECP256R1_SHA3256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp256r1_sha3256;

localparam int TEST_VECTORS_SECP256R1_SHA3256_NUM = 263;

ecdsa_vector_secp256r1_sha3256 test_vectors_secp256r1_sha3256 [] = '{
  '{1, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 264'h009364745a6a2d69f2283698fdfbee7b13de20bc93deb0230a9af3bd9fddf04401},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{2, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h8ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{3, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{93, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 280'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e0000, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=280b(35B), s=256b(32B)
  '{94, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 272'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e1500000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=272b(34B)
  '{98, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 280'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e0500, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=280b(35B), s=256b(32B)
  '{99, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 272'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e1500500},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=272b(34B)
  '{114, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 0, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=0b(0B), s=256b(32B)
  '{115, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=0b(0B)
  '{118, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h028ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{119, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h6e9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{120, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c3ee, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{121, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e1d0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{122, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c3, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{123, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 248'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e1},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=248b(31B)
  '{124, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 248'h9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=248b(31B)
  '{125, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 272'hff008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=272b(34B), s=256b(32B)
  '{126, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 264'hff6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{129, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=256b(32B)
  '{130, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{131, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h018ab9effc67388040d19b92d2e9fdea124fec6626e540f2b02edc15b83a73e8bf, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{132, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h8ab9effe6738803ed19b92d2e9fdea12d61e70cb9711b5a64768803241ad9e1d, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{133, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'hff7546100298c77fc02e646d2d160215ed6cfa9486c1d6abd4c4ddb50ac1ef3c92, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{134, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7546100198c77fc12e646d2d160215ed29e18f3468ee4a59b8977fcdbe5261e3, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{135, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'hfe7546100398c77fbf2e646d2d160215edb01399d91abf0d4fd123ea47c58c1741, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{136, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h018ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{137, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7546100298c77fc02e646d2d160215ed6cfa9486c1d6abd4c4ddb50ac1ef3c92, 256'h6c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{138, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 264'h016c9b8ba395d2960fd7c96702041184eb9bad38c76f7f19ff4c7fd7e61ad606a1},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{139, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 264'hff6c9b8ba595d2960dd7c96702041184ec21df436c214fdcf5650c4260220fbbff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{140, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 256'h9364745b6a2d69f1283698fdfbee7b142139c1e637988485a739f2dce18d1eb0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{141, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 264'hfe9364745c6a2d69f0283698fdfbee7b146452c7389080e600b3802819e529f95f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{142, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 264'h016c9b8ba495d2960ed7c96702041184ebdec63e19c8677b7a58c60d231e72e150},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{143, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ab9effd6738803fd19b92d2e9fdea1293056b793e29542b3b224af53e10c36e, 264'h009364745b6a2d69f1283698fdfbee7b142139c1e637988485a739f2dce18d1eb0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{144, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{148, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{149, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{150, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{151, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{154, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{158, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{159, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{160, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{161, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{164, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{168, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{169, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{170, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{171, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{174, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{175, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{176, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{177, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{178, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{179, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{180, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{181, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{184, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{185, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{186, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{187, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{188, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{189, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{190, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{191, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{194, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{195, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{196, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{197, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{198, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{199, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{200, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{201, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{204, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{205, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{206, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{207, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{208, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{209, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{210, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{211, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{214, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 8'h00},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{215, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{216, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 8'hff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{217, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{218, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{219, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{220, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{221, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{230, 1'b1, 256'h9bb676eec3b5bdfab3f802242da6ace3af94f785c4ab299df8b02a9f0f76ceeb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h64a1aab5000d0e804f3e2fc02bdee9be8ff312334e2ba16d11547c97711c898e, 256'h404a1a6da158ae1473fce08d338b8d6410a6a5903358b23fdd3a54fee2c2742b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{231, 1'b1, 256'h00000000713791d986ab76aa7cb5c46cf5a62351efb6c1cde74a8591d9c2fed9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00a9edb87925684bcc5b92d0f7455123656e3498a0d182be63e2e6077c2b43bc6e, 256'h2c729ea1b01d14ee8fe702096cddd9394e351d801411ec8eac6b758475ea0070},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{232, 1'b1, 256'h310000000051db6185687c0e1d43cf6f7302a7ecf3fe3d6bd30b5363dcc85614, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3fba20ca893dcaf04e89141337a96abc7e24e026a8ff4c86d950de1c31b64272, 256'h6be2eced4ce388ff8026dfd3b658144f30931b7083ee2af06e75158c15b12249},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{233, 1'b1, 256'h80e10000000005f3acf7efe73a0182b5f719824bfa118c4925a1e8e0f194add8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00c5aa31116f6006c479586ff7070014a35f22166701be8a5f1f1e9a43cb27dca0, 256'h68d1cee35ba3893b9cc3b5df5ac6afef55ebdb7ad9236b1fa8e438a538f8cb55},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{234, 1'b1, 256'ha4392c0000000005c4dc1e6e2994620d6a959373e62fa5f6e84cabd790d6e56b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5b5b4d890504f56c16a4ac7947ac0057cdf640d2c39bac09fedc648bb0a16f1d, 264'h00f9c12e73a56d799e2827538187f0ed0ec331f6f0c089a4f6249d04c1b0c5cc8d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{235, 1'b1, 256'hd7cf0d00000000000e615ec0f55109462536b34045963901b95960c6cf5296a6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4338e710478e8b922e50dc947f6fa0cd1903106cf02ee0742da69e8b624c5b67, 264'h0090c73bd0fcd07a4dd4a3664d559bd4795ac950d89463680852d33915de1a5745},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{236, 1'b1, 256'h8b9d7d14000000009051340f34c75a0e78f4a191b3f908bfdaa334f32eb47b51, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0fc97d7744e0b2762e6b48730d44c758ab238136a72693ff27339aaebefad581, 264'h00ab68ec80cf4afcca0f7d75f3c4b00e34ed4fe9101c98ed4d8c2f97eb865b1683},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{237, 1'b1, 256'h432701b4c5000000004e77e86a34ff07f3069a9b547da784a05d7d5d950984c6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00825f0b4230e30182b24b65151ec83d0aadc63ecfe0a91b5879ccf7fcce9eb40a, 256'h47f0211ad5471d055fe07c75f37f3fad8aeeff1ee11a54a17bab35212c46d5d6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{238, 1'b1, 256'hee4ea2312d5300000000f10e2378adc2459d7728a0eb1c3fa70bf25ffdfc2d9f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3fedd83579431889710b67b6454d43ea7eddaaa9da950424e2c4ac730065a822, 264'h00b50cef5a9da8323fccd5bf13260dea6517c8ae6ccd6495f9ed7494cfd5891573},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{239, 1'b1, 256'hb519e0108d975a00000000885c7dca69fda64d70ab959d0a99034d75dd180ce7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h69ba62b020a36333f7a0716577dd57d280132c540f66b9e2fe8d470121e0f135, 256'h66c7811587cb9247ec6d8c223b4c6d5533948fbabf072973d74cb19d3b2c91a6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{240, 1'b1, 256'h0ab9f26cae100d3f00000000d72de1818987a2554c6818367ae35f6d08dc2478, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008bb763097d8ca8e9cb84e111f361f47de93499f50bc85401ea96a61d54fad7a8, 256'h2587b81e277283d5c139b8e9a5f4aa0bb0b1c2b28963efddbf73a0eef341659a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{241, 1'b1, 256'h20069e1ea6d4dc3f640000000096664b82ba5b4b6bbef31881c2e21cb8b32bf1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008260a1eb8ba8b52db95b0722887920a1f9989dfa1efd420d1f8f9ab3df0cffce, 256'h6752c5687e6889e008eb9ad6e41933796b4adcd6018420fdef250998f6adf603},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{242, 1'b1, 256'h88c1ae896d5b1ee1e1280000000051e2c22d970dc99dcebfd57a35be0f5195bb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b809c133b30c3a8ff11ea9024b131664b51c2768afb8536744e041015da93806, 256'h6cd015a49e19b260da6cd32a94806fb8bdceec5dc5542a7b2b938cce75137f30},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{243, 1'b1, 256'ha8dd2ff8e9ecfade5537f2000000005f36a2ec63912dc97f1b148cca8d3e986c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2069244f8e72562406d631f647a141831aca5907fbff09932797d8305ad3c19d, 264'h00dfb7a3ae1a4bdf76987d7de404c5d8b7c51a6ae8dbece9de345a4b71cb5e1f38},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{244, 1'b1, 256'haf52ca1d210a9ea8ae35e8fc00000000cec8a7eb3b52686105536d8fc3757f7f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4d82e457954761001da6c5dd0fb45d3b8aae12a270cdc5b97d66f810e3065326, 256'h0cc6217e3aee3839fd809b207d47dea412991932adb2de18ee86431452c22595},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{245, 1'b1, 256'h913090d6f8bbd4e10e2ce1c5450000000016451243b9db301de24772cd781cb3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00a81c6258489e10bb1132a6f81f76c31d7465869708d89eb018c51bf774e8a093, 256'h304d75b7bebe9abda5daafc419a765ffb8e5c02dd91836c40c430f052d5ca59c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{246, 1'b1, 256'hc1cc5ad98460c3b9e3852479a3df00000000808b0b9e82f6ade0de221aaa7ab3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00e8da776984d6af2b8d523d1bd6fab8b25409e669d172ef51e104648c1bf0dad1, 256'h49b4170fed1cc59ab000087a2c091b3f69a66c8562ed350472e982bd31a0d09e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{247, 1'b1, 256'h777e0e4f4ac2bb3050202e89f5cb690000000030c36872c4a1b6f19c1a447203, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00c53d293775c5cfdb879b67ff4f4792942132c35c9dc7f8fda8b3a00967c75b47, 264'h00c36045151f70a5d6af2fd27cf1f13cb308b2e847151fa4b47e22f2df6220ae95},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{248, 1'b1, 256'h8b15a9990c7fe432804ea9a57b1c8db8000000000033521f6cd85d48845871b4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h300ee6fa4de853ac6680302a9c439b82dfd046c314d7bbacb2e01274e61e9b54, 256'h0bb2b62f11b789848648fab7e0c46ca7b09cded01887ef6bda9f871bc5cc609f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{249, 1'b1, 256'h2b623d836940fd3a612348a20a8d1caa00000000ad69c80f64d89f5f050714d2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ac58a18fa5973efb06adba842affbd256a1c624606b146dae5a6ef85992cb428, 256'h48b4ecb8697e4cd20e0f30721ad94f4c18943879ce5d99d8c000d90465138bd0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{250, 1'b1, 256'hbac4743859e5588409f25335619fe1c7d2000000000056aaa54240b186b1ebc1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6ebc2857fd53656b857005eb8f95c4f6fd3c99f9636a028e5244edc60bc9e18c, 256'h27719f12eb1de6cade547cb98523bdc7108622240f38d12f415c79cd0b1344d9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{251, 1'b1, 256'h7eabb2d7d21887903ffba869f353928bd5000000002d3e45954e4b6e21fd30d0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h67e8ca1907624419e3ccd88002dd7757f595abc84bd861cd0198364a4571ff6b, 256'h0db40b6a7200cdc1a09df432a5a763436ab4130cbdee024dea2a3ddd6c023ed9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{252, 1'b1, 256'h951cd3b90eec711648999d2ca3e8e821b86c00000000574333322ca94097a491, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00f4d8208eed5cb4bfe4ef6ddbbc3742e780e4212a39cf79c9f85605ee64a962cb, 256'h43dee8a3c45a45a91e83a18ff3f881047b4fd6ad3003b3af37fb8211eaf7d584},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{253, 1'b1, 256'h01ca3636d480cdce6ee63cbe3665c7bd88995f000000003f5d61628138af2b7a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3363ccc93e2413e47528ab086408bc0521be73353f2c2371bbf2d9dc16e63fb3, 256'h68f3d1074a2e06d33fc19a567a8af0edcae923560cf38da2dab82e2249c8dbbd},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{254, 1'b1, 256'he64458ff971279b567c8eb016ac86c39f963cbaa0000000056fbecb71ef3fd7b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h0084960758125ad8de3df0c113ff35f1644e4d43f661c2d81848f3fe4e55846f18, 256'h5983630fc8975bab570d2c9f3cbbdecb4dd6179ec497aff312d807ec26ca940a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{255, 1'b1, 256'hb15bafa66eaa8c73cedfc9568ac5a41a5b0a45e38e00000000f88ffd117bf4eb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h06ca924b5686a22f2e39c0f980fd58d62bbaf33c3a57f98a315332121e9ba60b, 256'h6516b98b31048722ca25e0a6c450461823c0a35f37d671439084fbc27c4779a1},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{256, 1'b1, 256'ha0daa5e1d6fb10cf91937045a9adcd668e53d8d302a8000000000223f8bb456a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0093c5ef07a7d955056b88cc8240060b4ffb42835a3df353cbe16ccb62eaf3f6, 256'h364dbea6d5ead4202d6fdc253bb0c2c0522b55823e8bb890235ab09ae9030ea2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{257, 1'b1, 256'h4b28f92a09aff0587c6eb0a61588a5f2d6b1e85955436500000000ecacd385fa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00835274f3157b737975486c73e5bbdd15b61e2ebb9e580911e45fc288214d2e67, 256'h1d5dcebfc6d3ae3826b9a3211f5e2249acc967eb47dfd41a849241ffe779154f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{258, 1'b1, 256'h1d29293e1f2113a0eec5780d25200ee18779ad86ca0431390000000088a9c6e0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3797916fb5c401a691b710050df3eec163383f855f93b61322a56d862ad5572d, 264'h00eb7bff4000738a83dd64082eff710d5eb619427198ac290b291f4599768959ca},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{259, 1'b1, 256'h3f466438a18ea4e57a572e3ee501d7919c87bb35179a13bc5a00000000023949, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h70992463694c845183db142a77bf5d73c17e9004a8b946b7b8eeb3fdf2b22e00, 256'h03843ec28e4c4d4f7726a5a5835575bb3e272f612246bc3aff288ac4a4e90c90},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{260, 1'b1, 256'haa2ef39293ec474361e7562735439b835b55d17b130df2421eb200000000fc40, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00aeaf228b41a1f311d4df74717f4134ee992e5f2922eec65ec83e2db82a866472, 264'h00f5ef65eb9fc3feaaac04f71a9a5ceb73e8cd6cb75b4595b39b250a50476cb68f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{261, 1'b1, 256'h1df7127ff896950a28abfee5f9dd0da5da0f5960cfb1d46fc1617800000000d9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b84dbbddd3b8a2ddf67d27e4ef886f72d90cbb7ec2d6883728b27842d61505cc, 256'h32be7f0ff420ae3be212beb4c276d93e2527b0964d643c5807c8ee711e66e8e5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{262, 1'b1, 256'h69e86af97404788bda6b6925dd727c578ada594a03d4975b545b70a800000000, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00f7f6782978f376caf9434941535e1c87ad09b9d39ee936145a0b53b9250fd182, 264'h00fb752930c84c29e49f81a997a4d0f00fcdcb4a2f2bf8049cca5d7cf70b079cea},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{263, 1'b1, 256'hfffffffffbda4755bba6de00c2701a0c6fd32c7e4aa1d876140f979cc80f34c6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00fb4b434112c1302ffd49ebd993cf5ec59729cbe78739db3c470264e378d56e8d, 256'h3aba99bd10be0fba04ca8d9601ae8f68ca7ffe5814f4cfbde78c1cc07a29fd8f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{264, 1'b1, 256'h22ffffffffacfab2fac775cbddf678eac83d9fa2dcaa8379ca3af3fb8dd614df, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00eafafe851aad76036013bd571772147b7257fb736ed7b4458e0dcf60a2c7b9c0, 264'h00b59c6409e51043b7e5c86a8d465978a4c8f78e13ef5b184fe5f46f201ff4efa8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{265, 1'b1, 256'ha92dffffffff4bf463c8eca0c62afb2c35c2a592ad8e8e688aa521a258f47338, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6c74d1679d871a46a43c3fe375e09d4f1b6413c59b5e070d7984dae0aadbc37e, 264'h00ff1d22228c9e9cf9958d677eed4c3a252b10273ce2d360457faabe7f7439c0e8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{266, 1'b1, 256'hd0fab1ffffffffbf5c5a0dc94820af6ed2c80b5411be656e273b963141464e36, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00cae28b592e2d5bf6f9ea541e70bceedd07adde40bc2b5f883d35ae9560fc85c2, 264'h0099eaffc16f570b7837d74177dae6e6cfd873ea89424581bc690d0e49c4218402},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{267, 1'b1, 256'hdf0ffccdffffffff58bc3fac8197329161b5dea9f0043e8cec2a9a631ea38cea, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6ce5133579dd044447206b9f6e1605d27f094b2c4466a5bf8e157873176baf3a, 264'h00bbe35524d9c1936bacecb6c270bf494eac75933caa8dbb2fef30f6572ed8667c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{268, 1'b1, 256'h4d77a2c899ffffffffb8c2d8566f592706ca04276262ff7cfdba0b2ad6e2a6c4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2855cf6e65812ea246e366ab961970d19387039a93f0bd406365d68b03566613, 256'h1b3a9593117380899d5c8f8f976ad4dee97db9f1225f735b1d41c2a115be93fb},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{269, 1'b1, 256'heef9d05b88a0ffffffff18a16611a3f3ac44331426f2bdbd5af203e092e61176, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h0090ed3aa89579b73477e3fcba9f52a5a64b9b6d83b475a3881bc0e63d74f6bf9c, 256'h04cb5e2ca1d413b37a71607d5b5fa72ccc87a2edcd5c7f30daaa94241b749920},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{270, 1'b1, 256'h7e6d3c190be6c8ffffffff27a4b129531bcb4fad150112ceeeeb8d10098dcfaa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h055e38188756831ced4b01e0f9d4db6b02293c7ee2c3fd47860d38377ee0f419, 264'h009c29f1688f16e111914d9c843c0a8f0306c1c4ddd5167cdd54338a4f4ab79a91},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{271, 1'b1, 256'h0edd238c04bee70affffffff0ae88780ec5271030a1847cd73f722925df9dd43, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h06b28cd8538d8cc563473cf6c7abb519e4c8bb4c37915ef76512f37de02c2164, 264'h00a62dc2afb01a1a9bc877edd54f25fd1f6d0378b3fbaa219ff9ef28c560cc8065},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{272, 1'b1, 256'h4dd115320049ee2e9dffffffff0de268e472eae1699ca5afb5c838313db94bed, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00c4b97652702efb1d1b67e966e88789efc0d9eb76d32efbeaf9c1bca36b2ea9a5, 256'h13e1b2358c7a34fef3ea738ef1a48fab63a2616455c81f8095394a2230c852e3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{273, 1'b1, 256'h1a1109052e9ab4f5dd2cffffffffb1e4604e058f3040a4af85f1f303bd3830cb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6a86100848566b5f5f89c13643515d81390952b6b5ce56b64fc3349e4edf21df, 264'h00c9ca4ba3a6fd501dae9917283a6851692f57dfbfa49d7a31aa937534df760c87},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{274, 1'b1, 256'h6162159e82cf80a70b34f2ffffffff193b3c777305a8fc809337cb13014edc7a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00c1ea204ee71a0502fc47de5d89fad98b897b5c308a4030b4a29de9cc39ff1704, 264'h00a5261798ed9665358c31a2368c6705b53b5d7d17023c365ae532573593934481},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{275, 1'b1, 256'hb35876d301bf4040fac24355ffffffff7fd82e02fe5885a42240d05fff5fc61b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b3c13e4907afa5a629398ff4fb50c48fae69dd3721a6f62ac13b901efcb4717c, 256'h6cb8a95728751b6274fb57e0e8fc87bd7911b1b94fb92edf09ef30fce410efe7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{276, 1'b1, 256'hc5ae766a399aa8c082a59a4f62ffffffffab6578abad5454b86f0be4e36bedc8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h009fafebd8841588e56116b2aa354557be814630bae5824e187405f3398f36bc5e, 264'h00f01264feb46aeefe68c967e439986f14aeb85ad99b520db572af8d1349d696a6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{277, 1'b1, 256'h619548e83b2bf592724b244359f9ffffffff7ed41c49517b65795ef980c30f19, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b45703f2c6e95c2f2378913cb78ecf7a01932b66d85e6f687dbb618b056851e8, 264'h00e1333352ea3ad42d7fd9a52a9b6dd1252848a180606d30012e142d135156720b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{278, 1'b1, 256'h2ca970c6acc18b4ad3b023ba01ac4bffffffff4fa0a25f4f35f9b408dd09517f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4138934da6329335702814333f4df8f907df7aa8e684cc38e2366961828ad937, 264'h00b90b1b0d77fa39c81f3df7a471499ebbe415a372e7c947eae8612646081aeb47},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{279, 1'b1, 256'hbd67ed69ca5085f9326153231b96b177ffffffffffb1a4447142406fbb23dd5c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00a52a6cca52d60aedc270cfd2fb0e0c2dde1ec4bb61434a7f11cd126ad46bec56, 256'h1dba92bb08e5665da3847abf695dbe18aeae37d9fdcd3617fab0c648f48d8ce6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{280, 1'b1, 256'hacfb85a5cfe484ca5801b819b3e4159dffffffffe10cb294343a640526d5faf1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b153363d48a58d339a7e53bfedddb63ea63484569bda2630d61c129a45d352e1, 256'h592dc8769b4834fae70f2cf3eea157ea9684c56d4875d296313cdf12e4939df8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{281, 1'b1, 256'h62c18f3f3271e3341a7d3033529b28a2c3ffffffff4e9cf2e8ef755e0953597f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3516e0c8c97110170a5121b5408043f33c6efbef0e5556165812713be6422ae8, 256'h5d80c5dffa87d3856083bf67beb27e90ebdc2e54d84760c1588f6432ca733195},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{282, 1'b1, 256'h2df78ec6d8628aeba725a007584b63636883ffffffff0ca2480cb4e3523b2daa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00903d8397244bfc99f2a677507db419597fef6f0cbfd49e0c022709c06c93e358, 264'h00f1705f4a19ab86893e0e022bca9081022764bd986c1c891eb80202ec46f50870},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{283, 1'b1, 256'h07fc58409c7cb5c7169a63d09e4de5120132b8ffffffff1f95f5e389535720ac, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3ba4d01ac8cbfc4abf848253d060a4e3faede188fd01c21657c20b61d1943f43, 264'h00ca3b5365ffbb98a5539cbe3e71b3d9fc59b5f1d5bee1122870e153ded9e1ce67},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{284, 1'b1, 256'h383dfba6e0aa10f820e15e27374c2eb6996baf43ffffffff66a94ff532236f85, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h741b76d33821c8cac2361048f10d28060f43e2c30b42b3f1b64a432f322e705c, 256'h37331cdebe152ff84bf909183069f278f8b0779042d5486b2d9826b42546952d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{285, 1'b1, 256'hc41a8affa1bbbe99587538b31e0b61f8b56ebe58d7ffffffff45e1ee3efb6c66, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00d7988135fd211a2cc09a4588f2d91de3a9a9498d5c5c3ef7e78e9bd80906a63f, 256'h25de3162aefbd6afedf01116b4e69d498eaefbf29599a7e0ab60614d64fb3db7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{286, 1'b1, 256'h26fa9d690a2129917bc3520b913f913f1f081bea9aa3ffffffff0fd642c24a4a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h14580cf3aae5ebbb74fed09ff193f347f69ac5b38435eeb7c38a0fd95f5b7ad8, 264'h00fcd923fdbdcecb3ece3bd0069c81396b4acf6328648fbe5324ae0c5a276fd87c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{287, 1'b1, 256'hb291bf1a8c66adc9def9a0a96da478aa1d09e06797adcdffffffff8fb0460842, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h130821bb00d0f4416ef06761aa283d35383cc2d46ad6be76c96d839adce2dbb6, 264'h00d9deef38e7d0f136cc535f1f8931f271cbf0b0d9e4e20fc8db7a1fb3c616bb68},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{288, 1'b1, 256'h81d64896fa11ee94e49755c0180cc0478de87bf9969ae759ffffffffb4b7f4f5, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ab4991cad903fc45f6afe22b939640736aec9788b9d8f94109343649d6327695, 264'h00ab126decd1743caf4b461a9c8029cf1230a54a0180e5225a79c075167c2911bc},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{289, 1'b1, 256'h3b88244a6ae111bc752afc8f997cc9ed1f9d4079a0f644f3d8ffffffffa41c42, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dc3b756b20b906f02dc03b46bbef56708be649bb4b23a41ac4333cd79d72749d, 256'h309dfe0623034d6441332aebb327bf5b0fb2f3d6df5a6c02d836fc908e37b0e0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{290, 1'b1, 256'hbae669421b6378571d97fee160d401bf8f4698bcfa6788a85be7ffffffff6844, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00d733b4391a4876d30acdb95977e4fdfded201e698e42be54c5c690b4c83c9036, 264'h00f55565475dc58e468b4aaee60eda224770c5b30517944c065758cd5155ae1251},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{291, 1'b1, 256'h1f52ed3bbbeeaa23026b261a17bc00058f2e37cba29772831b7ed9ffffffff02, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00aa9ea086e301728e0cac7568bf64095b9f51d070edb46679a9983500245e3468, 256'h3aeb2415f10625c3a4e818da7ddecea27f56f0a393920f6a5d2f4f3054e2131f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{292, 1'b1, 256'habacfdf5c9518bfcd685890b4e11728fe6bb738a9517baacd701149affffffff, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00d5a6ffddece918c5fe4e7d3a11344612bfb0cd2735ce071dfade01244c3b303c, 256'h0ff4ee3a70b9984e49277b3b15252c9f255b9ed51c7a4473cf55a7955083a985},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{293, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h58e71ffbfd2eabf4e4a465f68100f3d23d4702537dfcca5ee89d18a75ad7f756, 256'h16535d3b19f050e443bf5dc38f7f7cda9df3798d4a2f65a413a9af5df002828c, 128'h4319055358e8617b0c46353d039cdaab, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=128b(16B), s=264b(33B)
  '{294, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h58e71ffbfd2eabf4e4a465f68100f3d23d4702537dfcca5ee89d18a75ad7f756, 256'h16535d3b19f050e443bf5dc38f7f7cda9df3798d4a2f65a413a9af5df002828c, 264'h00ffffffff00000001000000000000000000000000fffffffffffffffffffffffc, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{295, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h0a78dad1701d0551089d3a0ee329a22a9d8bf4263c8a50e0668d24306cf0240b, 256'h03950b34bb638c683c167a00ac06232c2ef1718d3ed7ebcfc145a41031b04ee0, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254f, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{296, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e5b027e1f5daf6e52eca80e35be28651bf849ff3de70d2a34c0d782b5aaad685, 256'h3c8e2cff9b02c90bf4d7d49c7ff2a261d26aed7d4022b41392c85a857d434579, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00909135bdb6799286170f5ead2de4f6511453fe50914f3df2de54a36383df8dd4},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{297, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h24c5462bb7d1f1763ce28b3a9f851d86d7cb4c5f7c61ed9ed7d397f1a920ffc9, 264'h009460936b6919f88646844b27503555262ef8a81e6704f43e07deda12aa06f4ae, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h27b4577ca009376f71303fd5dd227dcef5deb773ad5f5a84360644669ca249a5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{298, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6226bb83d3cef01ae27b7d04a905397682d5e4a5964b5160dba8a055a2e2aeca, 256'h7a3630d49d999d0e85e59fe762c9c567cb767ca2a0a7a7756ac917e6085b18e1, 8'h05, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{299, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h65af8c23310fe060a09e7366d82ea35f48f8e2c682eab3783de7d9711f5923be, 264'h00bebabfaf084741fc806b9698ef87c9459246b7846fa17400094ad0bb222c2cb6, 8'h05, 8'h03},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f26ea876edab91b4070c5ec6e36663fff86f1fe5ef73938b227766b1805773cd, 256'h07059506a5296d5766d4c55c06eebccf81c04e52cb14c3b198a18808d570d417, 8'h05, 8'h05},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h7811e16675799076c4f5ea78e5f833be4649925165672057443c436cf4017e0d, 264'h008e377d53fecdf1556b1cdfdd8270d920cf7c6d32c946af2db4c864faec6b1eba, 8'h05, 8'h06},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{302, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h7811e16675799076c4f5ea78e5f833be4649925165672057443c436cf4017e0d, 264'h008e377d53fecdf1556b1cdfdd8270d920cf7c6d32c946af2db4c864faec6b1eba, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632556, 8'h06},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{303, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h03c840f0fcdfbe9cba931726d54a1f9553732be832d8ab701aebade4524b736d, 264'h00942379f10b74b70ec5a06d31c7b65eca6f77a047e25736aace32cf46edf9e90b, 8'h05, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc75fbd8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{304, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h4b2475ae911ab3e3334bd5acefce2225e35ad7f4523df52c13f581b87898cca1, 264'h0095575d5296d1bd97efaa74a12cc0df3d556a614f176c25b06348af8d304ea6c7, 16'h0100, 264'h008f1e3c7862c58b16bb76eddbb76eddbb516af4f63f2d74d76e0d28c9bb75ea88},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=16b(2B), s=264b(33B)
  '{305, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h211cc26f1f60998bccfc6ae65cfe8f1bf2e70fc28b5aaf8e2a297f3f4460662c, 256'h3ffc8dbd9b58a341d5160ff03b7a503649967a9a937edbbfc4bf154aa6e1a0ae, 56'h2d9b4d347952d6, 264'h00ef3043e7329581dbb3974497710ab11505ee1c87ff907beebadd195a0ffe6d7a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=56b(7B), s=264b(33B)
  '{306, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h0a7bb520f0cc16284831167d3622b276487a7bbf41bf911d367b484f1bd81a0c, 256'h0c30d573d27d44e68fb9a109ac7faad2c57ae09de30d8203ab409cd3ca63af3a, 104'h1033e67e37b32b445580bf4eff, 264'h008b748b74000000008b748b748b748b7466e769ad4a16d3dcd87129b8e91d1b4d},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=104b(13B), s=264b(33B)
  '{307, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d528a48fb391dd490d3f32810570613d16fe2709b82245027705e359549b0e15, 256'h5f4a5ac279d55c9ea6371f56403f816ee723632911df9804f01c7fa289eb2361, 16'h0100, 264'h00ef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=16b(2B), s=264b(33B)
  '{308, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d1f035f0a28c0c49e6248ff373874da5b26b47e7cd89c1b3bd15402dc9bd7b62, 256'h7a182a1884f30222976579d766da681a7f31fe55b14e770dd0f3f1c09654b29c, 104'h062522bbd3ecbe7c39e93e7c25, 264'h00ef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=104b(13B), s=264b(33B)
  '{309, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h07df495050dcb1738f4e2aac5ba2c8a1f8e09d262a3b001865af3fba086d7aa1, 264'h00b596cde482a6bfdc5e49e4069fce7c2d1145d1e0f7fed63f9e848446fae479ed, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc6324d5, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{310, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00ccd70d8730532b28c78c27dbd3043fdde3e96f10ede406582c9cba2618dc03c1, 264'h0095d592c366bd189683fd581dde22fb91176b55d94e48dd81467234777d8c223a, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{311, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00ccd70d8730532b28c78c27dbd3043fdde3e96f10ede406582c9cba2618dc03c1, 264'h0095d592c366bd189683fd581dde22fb91176b55d94e48dd81467234777d8c223a, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{312, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00fc13b37baba182ba13dfc8ca74f5896483378aa9bd6f0aa931877ddc5e77262f, 256'h1bf8b9cfdcbbe0d62eed81e5874310bd51178d1c6d01b6929a345d94190fdf3b, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{313, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h20adbb6cb9e09ce8ee4b6bdbc2e8047a0b9dc811eb415a2a258906efbd8a88ce, 264'h00c16b2111b5991d98dc4c935da619b55f784c79f000830d514ffeb6ad3fcf0640, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{314, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f033aa211cf11ee61c247567974fb8667c78f13a35bc2e6bead4436c261f144d, 264'h0099b4d07b6ce8008fecf8a4c4af561b972b00e63443a2f20038ee84ed0c238a3c, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{315, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00bef2538da3d07158791556b2d0297ca9c1b306459c9323ce7d07a21282de1ace, 256'h4e400c8e4eb57751faa0dde6bbebf96faaac9efc80e3de768fb4f5a37f95ead7, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{316, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00bf2570b58f38183fabca3ca72255bd4651cbb7e8292287809bd8e5c285d24a53, 256'h2f859b7f75c2f5e8d3791a5ccb60fa3888895c63237c9ea65e43f87523e104e5, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 264'h00a8ce483a42fb3462047c96ca00d1ab83ca565b2724cca9ac14411dcb8ee7e803},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{317, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h009ba8f147332270987e5baab2ab0a4ebc9968eb8682c2872266a22b43c2cf55f7, 256'h728d552fc65b5a3c7cee18876f1d8b46ae60153aec3b8a2b2c2527979f4a7d29, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{318, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d9e64db2ea560162dad3ec67d6ebaab9e821a81da8d4584f00fb14813c7e96e1, 256'h53e9e96e17eb05228ff3c9cbc5318bbb87e88bec489dec2be7a20adce06cf8bd, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 264'h00aaaaaaaa00000000aaaaaaaaaaaaaaaa7def51c91a0fbf034d26872ca84218e1},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{319, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00857c58d9010d1f8386e279cdcc369b32a8960259a3a646f6d89ad5273252f3fc, 256'h65d2384cabf6a2158b1cd1b2e2477d10b1b719125e9226e99ae90a7afaab499e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h1d109296e9ac43dfa92bcdbcaa64c6d3fb858a822b6e519d9fd2e45279d3bf1a},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{320, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h0089d887b0645d2f96b407b080cf6db3685cc9d4454d35a5ac7983bb5ebbfd2e20, 264'h00de4fcd410c3b6e11f5e4cccb19327c181c43c2d216869309f22495d34ee2796f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h027d377d04715e43754629961c6233961b921b3283c33fcb541cc27285092e8d},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{321, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h040924291aa7975fd04f8b2e923a1f9121836fdfbf2fea123cc1870f4f6cc0f2, 264'h00c510ee34a325e772d232b576052f96d3ec4a33b086508682fc53099c0cd48e45, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00ce1602ee5a6d686c5b8d8a3f44f419aa6064f0d35323341d77a65a4bc9e1989b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{322, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h3e7ed2fbb89f7b643d4ab44895ff9fb16e8be7a8649e4ac4ee2f59ec8f68fc63, 256'h4ca91cc26043a8242e2969c871d3ca9833148135b27d377198182ceaa7e70fd4, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h328ab273ff681a79a9662dc174ee014ef73d597d32ef42b17f443a33f5e430fe},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{323, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e67f559f552772b174d377b239e60750299d379b6bec6fc93adf040269d58c42, 256'h6c397f7984a149f07bf79fbba3b18c925a797cc6678e2eeabec47fb4ac461041, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00ab27431e81a7976e62dc174ee014f0479c909f17919ec453013b47f1aa221858},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{324, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h0088b1d30e29fe0edeb93ab469d2698d0fbc2977f77f48293d0e87acc0856a51fc, 256'h3d1b4f23fa3f6ef26f0e94cb7a63907b1923e30d08197115050b9da98a2b5f56, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h564e863e034f2edbc5b82e9dc029e08f7c3a43817c25ea210ebcc52057e10b5f},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{325, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h23a6ed2b1064923104d08ee4392b44bb51555a395477dc52546af6c787cc65aa, 264'h0081105b8c72c357d75215b210286df781d6731c4f0b87e9fe7066489653dc35d3, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h31f2cced76db7b4d74ee014f047c96c9f3ba3e21f11248bcf451526ac376c54c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{326, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h592d27cd81fbb61ebbdd782eaa1d86d53b59eaef43496677c345adc9896c562e, 256'h355b8ffda4f8683da98653f0d6067bd8134c5c3e22e3dcdee6a5cdbd826f4915, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h668fcfbedd4eed7eb6840c7f6cf1e3dde504afe5732ee0e1bcbeee15b94a2c64},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{327, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h008c4aa42ef47c4e2d7b60ca2b5a0b3038a9f8e7ee1de77d299286db3cd635b754, 264'h00f65438558a2271c9444b77405a1f97e84036c3146c425006e65be83f97e41191, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h637e57bd4f085f9d3be20506bbc2b8eab268a33871b19da56b1ba0ac25927bd1},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{328, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f5618fb978b70f15b8e07a74edfbcea775dcb92055f9431b816cd4cb5d4fd63c, 264'h00bd1759fd35bae79bf5bb0394646b14fbcb1ed2614fdcc9a9f53663e09f8c6a09, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00b0a105281711f1755bbfc1a0b6ea67add1085e84b73016989e20a90be3504d22},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{329, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h53c143435247e1e2144c4c32cb1c900b8e9cb160976bdcda1b24877ce7266a74, 256'h41a21780d91554d349a4c7c61f799bda9ddc81a66323078245dcb3960417a660, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00f177b6b38b29de112b6a1921aacd9c95bf24356c916075b623d05899bf7945c4},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{330, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h0093486f6653c2906152eb9d1c2b28e51c085f20ac54016a808f6e3c6b2cdcc02a, 256'h35439b7b9ab9e86df0ca617737b49f28badf8f5636c9bbaa199bdd20063ec7ff, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00e2ef6d681653bc2156d43243559b392bc161702b7ba94ce753e6e670828f6637},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{331, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h5f2e06f0ec92b6499eb7d249ff0147639253e7abe0e4497226336a5c94caa777, 256'h4eb3c28acf5012ba023971416c600a10fb6d28a23f3a2c1f77fb0686d06cdf80, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00d467241ca17d9a31823e4b650068d5c1c39eaaea65f2241883fd744745a586aa},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{332, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00c2af0b9da06d54b1a5ff93800b579cbce295d0b2719da307b028bee3c657424b, 256'h28c4928f185f68312b47de31ad87fac134de90cf114cc85d45a8fefd9a3a2350, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00e70b0176ad36b436adc6c51fa27a0cd50ea5f5c07d1d695135b0128763225ef6},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{333, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2a3c0253d54dc8a2a72a31f815b0bb6c36d852f8db14edf1e1b71cd3a7389a49, 256'h4891bafa1767b85e36f7507fa5eebd3da0024208fcfef28d56cd49a980ba1465, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffffaaaaaaaaffffffffffffffffe9a2538f37b28a2c513dee40fecbb71a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{334, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h3dd345114090328ccc0bdeaf8269396593645720b0b326849d1fe81ec956f996, 264'h00ceee0a81d7f65e1205bb1b6963a8e0facfd2a6124701b1a152094d037a216f4e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00b62f26b5f2a2b26f6de86d42ad8a13da3ab3cccd0459b201de009e526adf21f2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{335, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00fc8207ca84c4af4229139de953da3bdebf694537c15406e172d631e98591f40c, 256'h34a0d957e39e9686914e98ea467972cedec5a5c6bb55bec7916dc71f7a4c6f77, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bb1d9ac949dd748cd02bbbe749bd351cd57b38bb61403d700686aa7b4c90851e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{336, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h60bf7beb808286d8abff60c20faed73997395124542e6b7672089d88c14bbed5, 256'h7f4af9606f9be0199e4145698a62ad2545123a49eb14e0c33317f6909e3915b5, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h66755a00638cdaec1c732513ca0234ece52545dac11f816e818f725b4f60aaf2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{337, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2dcd699362d3665b6c9260608b3faf989d45ac15b9da41fb348d5520ecdf4e04, 256'h03e483670aadef4615c7a13fe1bf3bf927b4e47a667660b505ba47affee92ab6, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h55a00c9fcdaebb6032513ca0234ecfffe98ebe492fdf02e48ca48e982beb3669},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{338, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e6205f87fa837c474a2badac671578de77d6a077cd286aed45403508767114ff, 264'h00c18daaf2463dea80300c1f4d7e25b9f603eefb2e2cbf012f31a819c91cad7cf2, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00ab40193f9b5d76c064a27940469d9fffd31d7c925fbe05c919491d3057d66cd2},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{339, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h357e7687a79243d5e030eb120a3652c2fb95fcb148813f3da95d044bdc31c8d5, 264'h00e3ed90ea73567cb36c0fccd021da4ccccffe40dfe1b603428969788bed4416db, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00ca0234ebb5fdcb13ca0234ecffffffffcb0dadbbc7f549f8a26b4408d0dc8600},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{340, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h3d9723a8ea5ebaffacab8bf87b1d63e42da7bdf94e6c2520a0786b7b534dacf3, 256'h3725db2fb27248274ac2e6212f9071495c90ae684d056b57ad18e72bce8f36b0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bfffffff3ea3677e082b9310572620ae19933a9e65b285598711c77298815ad3},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{341, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h4bab5b68667090ed13e5658cfe68f1247031aee80a8ccb52ba0505752f7cd3f0, 264'h0085c70129c1715d9610a41bf7a063b81c1bc7ec34bb6a1c95ccd08e09f1476343, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h266666663bbbbbbbe6666666666666665b37902e023fab7c8f055d86e5cc41f4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{342, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h7801780aaab4aaf31b7c94069609a5ecf623a6dd7e97964061c6b3e4103bb84a, 256'h59c111796624cccbba09394bca04af79a31cbd36176d2ec4ceaa700730d57300, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bfffffff36db6db7a492492492492492146c573f4c6dfc8d08a443e258970b09},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{343, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h55b0451d911e9c64516ac9e9da3da1703eaaa46a8b0a7025c8c5ed38b5474713, 264'h00f1fde0cdee830bf169da9ca3d70d56f4607989873fbdcfcbb740e9a42faf860a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bfffffff2aaaaaab7fffffffffffffffc815d0e60b3e596ecb1ad3a27cfd49c4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{344, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2e19ea3a973a4c155814f8a7b641e12477d288f958b74f6031326356f5061fa4, 256'h1acdd1be10c052eaeb9c22d3f04cfec6e91bd23d6d3996eca9cd485e50e85909, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffff55555555ffffffffffffffffd344a71e6f651458a27bdc81fd976e37},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{345, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6eafbcb683e05e0bdb2aa0ac0686f60b34ce66761b7ecffccd3da8fe8799d624, 256'h4547b4aeca8a8e56dba45750cd9fc4f0e3f1333dcb855566c29bd14457cf489b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h3fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192aa},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{346, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h50f51ce959e24ac86b1054ea016c57d1da5f4cee008dd800757a817606234f78, 264'h00aa17f3ef6f7a6c51381c63d66697b1b5c196eb1da73d7b73c33f9115d7432d23, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5d8ecd64a4eeba466815ddf3a4de9a8e6abd9c5db0a01eb80343553da648428f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{347, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h009c8ef36f19815572db154e8f47a8dc5cc807d551a7141fed8a2c15460fe7ee10, 256'h660b936644e1ccad24578811dd45a325214e28a78e99a0ed2df7354fe9bca0ad, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 256'h56be8aaebb8627ef5e37057feb3448f726fb605312992466ee8d9ed7cd43c1b1},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{348, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h009c8ef36f19815572db154e8f47a8dc5cc807d551a7141fed8a2c15460fe7ee10, 264'h0099f46c98bb1e3353dba877ee22ba5cdadeb1d75971665f12d208cab016435f52, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 256'h56be8aaebb8627ef5e37057feb3448f726fb605312992466ee8d9ed7cd43c1b1},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{349, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f2a3ebc44fe94406cd6dc9bfc79a84600ae568cf533131e01505012649e39b8f, 256'h0f886d549f83aa61ecd1eeb77ba7256e984f088c3b9183e84a16e96f93860e4f, 8'h01, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=256b(32B)
  '{350, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e30751018c302c6916c21e2239baa41f0e69c5acfc371bb3e376ad364ea63802, 256'h659cceeae0cabfee3ed33abacbc490e8716b5fbf11137647b524e4b855d7d659, 264'h010000000000000000000000000000000000000000000000000000000000000000, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{351, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00ef28340fb027dabc05a2bd3be99c6cc2730ab0c3d8289e6a242f2b76cfccf9a2, 256'h405cd0530183db6640119a20ad9c1c24ec87d4d9d5de42bffab54fd6cb6f9ed6, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{352, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h01b4e8eb0cf6f321006fc107246c1996f7034f56d82706cd8f14f05da0a7c514, 264'h00f158ad7ff3c6a08b2f057c6c28255f9513811f20ab18f7104df554d591913f78, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{353, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h0b1cc580bb6f71e4bffb731a1e74f929c04a10ff94ac2312359d3f13213c3b4c, 264'h00870213c2ad3665a3d243dcb55780e21c8601c5f9803f27e31ff22f8ce77e739e, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 264'h00b6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{354, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2699736fdb603e90b1d9a04fcd90ed39756ed567214033ddb5ad579213089d2e, 264'h0096acfb0baeec9cfe2df150aa06b01ba58d03162b497c57a0d305adb4c5f7f375, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 264'h00cccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{355, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2a3021069e8841f9d69ad4c2992b02dc7a2f5447afa55a4683c6451cdc4e7286, 256'h00ca4123520611085cb10ea80bdb851a0b09dd79703c420606ff658dba94c345, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{356, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h535212040d83b1802cd4a9c0b6ceb0a89de68b794ddf979c2ffb9a72e59eea00, 256'h7650166217eb39f4e03fecd48e9e7448032da261caa68d21df639ba68ee667a6, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{357, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00884a86a89981e216732916569f9e3f203806359ef9b9ced61ebb82d5f8030045, 256'h079ceef71b8f9e1deb29aeddaf3bcc780dff88f92b705c68f572ec481139b84a, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{358, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00cdb031f0e0bc432f0b959bc270456f6a500635732c76764010a5ea20f54a71d8, 256'h5cf6ce18411cdcb5056e4280e449c3ad6df90f9ae2dea4abc08280d99749643d, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{359, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6309ffd3c559fe1b0967213461d884b58d1cd549dbc297101d9db5a7e3fcf3d3, 264'h0088f5fa86bd31043ca6077cd1da4b283f4179a23e9d680f66a2081ac502732714, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{360, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6e564ff8412e92f5ee23fd299c92c57eb6ef0cbd17c28721b92625938d0eab1c, 264'h00ff8941068815c9ad2d3b7f05845c41c4acebb92b3dc155aa7a51046948a4eed0, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00cccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{361, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h0083fe782d906023da7ba700d097f8cc9618cb23f1cd89c213b98b8f9ae8fc023d, 264'h00b15de38b856db24d4d6cc79b6d761fbd9ac94dad5f172883ba09278ba86d9955, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{362, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d1dddc947aaf9e6930cc46072f2cf2b68eb5e32dcf4ee84ea0647a201b299fbc, 256'h6b382061309943abefa5938e8465e2f6afd051eab974d261797cd483934097a4, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{363, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d17c1c5505bc710145ef74984864fe861e64302c16bb4a4bc69b47507b3f0235, 256'h41480e047b19bfe4bb885ec127cf254db1041ae1d5e8fd77e08294d398b62eb0, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{364, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{365, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 264'h00a8ce483a42fb3462047c96ca00d1ab83ca565b2724cca9ac14411dcb8ee7e803, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{366, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{367, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 264'h00a8ce483a42fb3462047c96ca00d1ab83ca565b2724cca9ac14411dcb8ee7e803, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{368, 1'b1, 256'ha7ffc6f8bf1ed76651c14756a061d662f580ff4de43b49fa82d80a4b80f8434a, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h63f01899b4b0bfe9dc9929fd4526919b981acda781044ee3d2c337bf5fc74830, 256'h591381bdf1b1a9b01020b87314a128d06e4833342bf232779f61480739613927},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{369, 1'b1, 256'h5a7a8ec92299354caa012069a923d56d0043b22408fb36ff8cd0ecba3aacb0a4, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h10228beaf773caeff22a94602e9eff1923dcc51b277f64b482ea63218c350b0d, 256'h2104c8343f8970a28c9eb221a63c857ef385e758eaccc5f7d2ae975553a1534b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{370, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 264'h00e6e1b8c20e9d00f0b6cf1b2c39cacd9c50ee3f990553250f074a4a3eed3afe43, 256'h52f3be1ae2d2f9b2bfea8e8c22d95af4574581a9f4b09a89f7b6a4ad1c5b2776},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{371, 1'b1, 256'hf3683c9e3da9a7f90397767215345efe3be07565f14ab80d102f50644b98fbfa, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h20f6203e48fc4c66ae8a74ec61d5124772daad058a74b871914d37dfe9d409c1, 264'h008b68de7a4786e29b3a726ea7fd8ef2a585b5c8dadf11281f2caa228eb3df3f96},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{372, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h207db605e42c96035d54352c5bc55cf27d5ded42cb6b42bdaee499ea64784db6, 256'h7f83c09192aa04ce038e861699a0f27ca55bf32741dbc95bbf997dee57f538fc},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{373, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h67c259a2580089ed52780755c75ea8a26b9057cc1995e4b044c8176cefe3cc7b, 264'h00d48f63d31333054bbd7fab676d207bbdc4dea1cf1b4f71aceb037b8dc7f79555},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{374, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h5dc675a2beae6deeb1ef682e922c5fe47156e069acd08073a0f8d9184d6baa6c, 264'h00e33cad4ce48f22ff6e50b47ba5dd44046a78ed7873cfd3a2c8b2d4b49aad2580},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{375, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h1a3b5c4b4a2fb0c2f9efb028a9efc78993f3151683cedf76214009ea418d3e5d, 264'h00e82e87332e7bd004cad9b13857939c01467fc1c3e4207efa45ef827985a82435},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{376, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 264'h008c44ef660ab8936fe01571168435c1918d005bd24ec76f72cea8f0faeb9f777a, 264'h00d793dcb3a6d47e2451e7d62e1c284ae25bbfaa0820f58adab79c201ba8d34a3e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{377, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h4227a3dbff7ac5353cd32c8b3456397a7ee7c0e6809615fcee466b1dcde3eb49, 256'h22ea6ad811b27f944abe70b47f490d255760f8c3562e6f7e2c1da3dbe45eb540},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{378, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h36636162db85e8d300ee45c51b9da00a7c2cffd9a6fb200761a647ccbf5d7e8e, 264'h009d18374cf1f87a9051e563838e75728d3f2ff7a86c10292851b6ce885c5b0c76},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{379, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 264'h00a637fc972f3800705b8d5293096382d1c1ae7f670be45011b8bd29059f3049bd, 264'h009c4abb6bbe06552d5d598b07728ccaed1738eac9fc985fd786fbc0a7347da828},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{380, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h76bfc74f3b488b34835aee96ee96067f53da021cff4020a10996d6933a27c032, 256'h2fd1658fe4e09b2e711b10117f5c37d9c3ea8b6f55cdf1e5a5ddae2c966d7e4e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{381, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 264'h008e0c35240e9e5b7bf2ab351afb13ac2655653baeabc247cab2c71cc40da44c00, 256'h079cbf8c9ba9b53608b219d6989875d960bdefcde224cf7ac6f8e791adaa4364},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{382, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 264'h00f6ceb6c8f76c337f51f4ec3859eb16caec969fc02a61dec1a70fa4223bdfb254, 256'h10c0334298a98a6e5c12e9c0cad587dcab43199b43cdf3785bd9c36b30925ccf},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{383, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'h083000a8e6121939f4b83612727b2091d8abbbdf9c92bf9bdcace8366150ce6f, 264'h00ba693f4e0b96dcbeeaa78c0d744365761151740323c346a54d74b332568d939f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{384, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 264'h008a1bd6ef283948184b5a32d31860e97cc0c450931f024c30bb3b261f2552cdc7, 264'h00b7e50c0513a8ec730d112109e92761a21151e4bec68268e5c79ef804b757deaa},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{385, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h0c18337b701b6000d3ce3574664c5dc44ead6a1f2ee0c27a728ea0b0f37990b9, 264'h00c31db9b199b3e1709c44a44118d1d7cb75324ee82ada2318744eb89651e6f6c0},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{386, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h2133d6fc78b394d4c34e173120b1e48c7fed7b89a03e55cab90b1367155b438a, 264'h009293e67ff4b981e50c48b0304f7b1e6b530416ee35188302b1dd2f21e5cb479a},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{387, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h3604a98e926b2f9d7585e341a5ecc73a4e811c5c8da82b65790ff8a117a75bda, 264'h00a0ff07774c9a0d4bf83db294b970f2696cc29a73637aa454d4d3b45eb964bb88},  // lens: hash=256b(32B), x=232b(29B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{388, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h6bf7e8f8bc3a5a2e2249c92725cf0dffa9b72ead3cc56d05107a4d587563beb4, 264'h00a05332b5b424d97bfc080fe0353470610931cd538d2e4bcf78c6fc59b481d271},  // lens: hash=256b(32B), x=232b(29B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{389, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 264'h0097e099c73088fc37052180d0483987e50c155c993cba2e6c93dd9bea5798e2c3, 256'h4a9ec5f05739efb4ea93790ea22c3fc423d0aeb109cd13fb1b44d87ea52ca71f},  // lens: hash=256b(32B), x=232b(29B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{390, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h3988bce3195aaf7c9b008a9f1663a5e13a8bee7ddba33a1bc5d55aa49fd3903d, 264'h00c39f614828e2f71a4c66d86d1c3ec7e283f768033cff5ed09e93e3218d9df1c9},  // lens: hash=256b(32B), x=264b(33B), y=224b(28B), r=256b(32B), s=264b(33B)
  '{391, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 264'h00c3eb2e8f78a31f221d6003b949f8df6c7ec1e0c53803231e12438cb2b1b1d9ba, 264'h00b97cc1fcce1d8ddbb5e1bfa6d5300d7cac155494603c66f7eee8b8e9c9643431},  // lens: hash=256b(32B), x=264b(33B), y=224b(28B), r=264b(33B), s=264b(33B)
  '{392, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 264'h0089e0c23ccf61e68dc0cb9777f18b18c84b2b02b4360c79eaa40d46ebe7f3d9b1, 264'h00a5d0164e398764e7d12d696750fcb092211c22dfdd3941e59cd73bc48eb91496},  // lens: hash=256b(32B), x=264b(33B), y=224b(28B), r=264b(33B), s=264b(33B)
  '{393, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 264'h00bbc1bb4ffceb61a0dbe5a12d9638dc9f004e797cf72cdba8d879fdbcd84dec14, 256'h65a7c17d9a6892cf5455a1904fdd9b57ce2b41549b9b2ca5d7d182c305e9a202},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{394, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h2f093a33c69eeaf847e332b12bd0758be41dcf75d8131878f16e6f121cb3f4f1, 264'h0093c304df074aef8cc2c8cddeaffda67eb2428ea7d3a113d51363e178d8068f71},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{395, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 264'h00b686774db39201a9462b96842adbeea16ae6003789bb18214dab9e5a758bf6ef, 264'h00ffc6b396293b94c96fcb325fae127608ebfd118a46f715b49b918caafb602a34}  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
};
`endif
