`ifndef WYCHERPROOF_SECP256K1_SHA3256_SV
`define WYCHERPROOF_SECP256K1_SHA3256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp256k1_sha3256;

localparam int TEST_VECTORS_SECP256K1_SHA3256_NUM = 256;

ecdsa_vector_secp256k1_sha3256 test_vectors_secp256k1_sha3256 [] = '{
  '{1, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 264'h00bbdbc26e1099b2713ada34df9cfa8edaf905a4a6d2a1f449f05de03df8c2a696},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{2, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'heb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{3, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{93, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 280'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe2510000, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=280b(35B), s=256b(32B)
  '{94, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 272'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab0000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=272b(34B)
  '{98, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 280'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe2510500, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=280b(35B), s=256b(32B)
  '{99, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 272'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab0500},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=272b(34B)
  '{114, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 0, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=0b(0B), s=256b(32B)
  '{115, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 0},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=0b(0B)
  '{118, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h02eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{119, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'h46243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{120, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe2d1, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{121, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739a2b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{122, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe2, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{123, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 248'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=248b(31B)
  '{124, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 248'h243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=248b(31B)
  '{125, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 272'hff00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=272b(34B), s=256b(32B)
  '{126, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 264'hff44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{129, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=256b(32B)
  '{130, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{131, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h01eb044a2e719d94a33837717ce9bc5ff94062cf047015777244b442e323862392, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{132, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'heb044a2e719d94a33837717ce9bc5ffbcb051537118436fac50f85c98319a110, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{133, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hff14fbb5d18e626b5cc7c88e831643a0057a4c0de23f3328c97b1e1ba9acb01daf, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{134, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h14fbb5d18e626b5cc7c88e831643a00434faeac8ee7bc9053af07a367ce65ef0, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{135, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hfe14fbb5d18e626b5cc7c88e831643a006bf9d30fb8fea888dbb4bbd1cdc79dc6e, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{136, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h01eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{137, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h14fbb5d18e626b5cc7c88e831643a0057a4c0de23f3328c97b1e1ba9acb01daf, 256'h44243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{138, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 264'h0144243d91ef664d8ec525cb20630571227c5815268bef4c2d8f46dcdba7a9dbec},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{139, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 264'hff44243d91ef664d8ec525cb206305712506fa5b592d5e0bb60fa21fc2073d596a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{140, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 256'hbbdbc26e1099b2713ada34df9cfa8edc3e56c7c02359540e308b81b1288c6555},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{141, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 264'hfebbdbc26e1099b2713ada34df9cfa8edd83a7ead97410b3d270b9232458562414},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{142, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 264'h0144243d91ef664d8ec525cb2063057123c1a9383fdca6abf1cf747e4ed7739aab},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{143, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb044a2e719d94a33837717ce9bc5ffa85b3f21dc0ccd73684e1e456534fe251, 264'h00bbdbc26e1099b2713ada34df9cfa8edc3e56c7c02359540e308b81b1288c6555},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{144, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{148, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{149, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{150, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{151, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{154, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{158, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{159, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{160, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{161, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{164, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{168, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{169, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{170, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{171, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{174, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{175, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{176, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{177, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{178, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{179, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{180, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{181, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{184, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{185, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{186, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{187, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{188, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{189, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{190, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{191, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{194, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{195, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{196, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{197, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{198, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{199, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{200, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{201, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{204, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{205, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{206, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{207, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{208, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{209, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{210, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{211, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{214, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{215, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{216, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{217, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{218, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{219, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{220, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{221, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{230, 1'b1, 256'he2ffb90fce551452ae842aa8dd047af56bf0d0ec8d3d141e30b36023b7c5a837, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00dd1b7d09a7bd8218961034a39a87fecf5314f00c4d25eb58a07ac85e85eab516, 264'h00b98c5232f0100d55db14eb0fe9e943fb45d8f192bbdd38147850f4d950f16a91},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{231, 1'b1, 256'h00000000713791d986ab76aa7cb5c46cf5a62351efb6c1cde74a8591d9c2fed9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00840a6cd819f21a2a3c3be7461bf516f5191c32d059eea09699ac4132f7948819, 264'h0094c53906a1595cf9fe14831b5298b4e297219afb895c18a19f4508fa4f6e0394},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{232, 1'b1, 256'h310000000051db6185687c0e1d43cf6f7302a7ecf3fe3d6bd30b5363dcc85614, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5928b7eeb84242914d4d5b871feb3b0d789455e44a41e3b60e0e43856a4a7a39, 264'h00d650930d76eb2444713b63b501a8e8b39615784306f1f2fa90915066e4f60192},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{233, 1'b1, 256'h80e10000000005f3acf7efe73a0182b5f719824bfa118c4925a1e8e0f194add8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2ff05b06077811e7bf8a1b8804fa6bb7db793b0a8927745f5b543998dab306b3, 264'h00c9e7da07e2b2d28f169924bab22d90a107ca97f5022eac08d0a4577f30d89988},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{234, 1'b1, 256'ha4392c0000000005c4dc1e6e2994620d6a959373e62fa5f6e84cabd790d6e56b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h19c5e74fd3ab3847d1ba8ec6ff682b184ed2ae466622890deb4206385c31b0a5, 264'h00c959ebce99b3446aacee56eecdbae1898fc71a6bacb4464a6a4b0276821b32e7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{235, 1'b1, 256'hd7cf0d00000000000e615ec0f55109462536b34045963901b95960c6cf5296a6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h54bb584a67c79e19d3f9627cc1eadacce8075e3f5c03e45c807b46d505ca73ab, 264'h00ab37fbc790a0400debbbde06b9771b63732d79de6a56e87275a968e0d4aaefbf},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{236, 1'b1, 256'h8b9d7d14000000009051340f34c75a0e78f4a191b3f908bfdaa334f32eb47b51, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h699d4d68c233f44bf1d3f70001a9acac7be906e09ac440c8d16044364696b94d, 264'h009990c2cd8d7c6a227dce6a94900bc7b69a8ee6cf0ba062767c09d9e5b12e413c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{237, 1'b1, 256'h432701b4c5000000004e77e86a34ff07f3069a9b547da784a05d7d5d950984c6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e779c882a97701293daa1413f9fe49ab97bd8f742331461d0e3b93333c1db5bb, 264'h00ad3fd904ab463ec8bc7ff988c142acdbc5dd73d8dce919b458987c1f32ba3e9b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{238, 1'b1, 256'hee4ea2312d5300000000f10e2378adc2459d7728a0eb1c3fa70bf25ffdfc2d9f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d121d4639e90e4741919d9cb3888d69c46d6fdc84980b5ecc249fa01cae19be5, 264'h00ac0559aa580e535e401ea9e2710f067a375ec69dc49fba668d7a14d8bde42d0d},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{239, 1'b1, 256'hb519e0108d975a00000000885c7dca69fda64d70ab959d0a99034d75dd180ce7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00de04d387ddd0189ef2ec494594ed056675788d6cac25f9826e50fec66f47be6f, 264'h00a55cbc3e87809b4dcc634cea32fc23cf7ac70f71ef1731de41414c0a71891cb5},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{240, 1'b1, 256'h0ab9f26cae100d3f00000000d72de1818987a2554c6818367ae35f6d08dc2478, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5a8d2d504831a047c7277d9c13f7f456fd9569a311c5be93cbfa9a3122534ff3, 264'h00d0f9586630564236e9b133a7b53202b29d3a3caeb28f5d2360adfea238f41529},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{241, 1'b1, 256'h20069e1ea6d4dc3f640000000096664b82ba5b4b6bbef31881c2e21cb8b32bf1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0e2dc3e0b7c51be950c814b4cd74b8707753bc5a7543d6589ae1464c93227bf7, 264'h009cea04df1218bb7a0c851da9fef4069cfca9fc00ef08c37976adfc4ec7b5e2b2},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{242, 1'b1, 256'h88c1ae896d5b1ee1e1280000000051e2c22d970dc99dcebfd57a35be0f5195bb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0c93646c509040bac868258bf3f2d13d26e98993e8680f0da846c1712be95109, 264'h00c65386f8b0a12fef25791cd93a045140af9c24fe3d3d700e02d23b1ce2da05f3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{243, 1'b1, 256'ha8dd2ff8e9ecfade5537f2000000005f36a2ec63912dc97f1b148cca8d3e986c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009906860d728638f6a260e13495f2c6099838e5c2f94828f10caf2c58970d3bf8, 256'h4853235fd511b8db3956bd25b772fab54bad3867d1c637a9984016f785fdc6cf},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{244, 1'b1, 256'haf52ca1d210a9ea8ae35e8fc00000000cec8a7eb3b52686105536d8fc3757f7f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c6d609fc861a35134b4dc180a3b2a7b13ad8477358e80286f90499c58bd37dd3, 256'h0978e0b21055dcc81844d297d6bbecbd074f09717b46c695ae60799d564a1f9f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{245, 1'b1, 256'h913090d6f8bbd4e10e2ce1c5450000000016451243b9db301de24772cd781cb3, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1496fd7a5023faf78b0e1008b054f25c509d34713d4594cfabf24c1b2229643d, 264'h00f660ac1daa7700a55189d6710a373b350ea2446ae76fc8a3522df3e01a2bc2f1},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{246, 1'b1, 256'hc1cc5ad98460c3b9e3852479a3df00000000808b0b9e82f6ade0de221aaa7ab3, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h31007f0306f171eb56c9bc7f7c0cd7d776acd86be680f600d3729aedc03aa9ef, 256'h59f529aecb6c8e7469830daea5065e6da8c349688ab4fa0ebec364035a68e58a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{247, 1'b1, 256'h777e0e4f4ac2bb3050202e89f5cb690000000030c36872c4a1b6f19c1a447203, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fbe1a139e3c74cef01d21d9c5a47a783080dbd9b86a202e933872a71a4b53838, 264'h00fe3164ad51c080ddd4126f42979e6b519075b2ec96060e02f9dd6fb6f9f3bfdf},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{248, 1'b1, 256'h8b15a9990c7fe432804ea9a57b1c8db8000000000033521f6cd85d48845871b4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h04518c6be6586ceb5559014ff40311fe7e6d0ffcdfc655b6a06bbe203a185ed6, 256'h1e0b927e43125aa196329bb0f09bf75d0481dba924f91e3e39e3e0878a972a83},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{249, 1'b1, 256'h2b623d836940fd3a612348a20a8d1caa00000000ad69c80f64d89f5f050714d2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ad67c0270ea088a9daa805788b6aa5161c6e7e12d237515518914ab66d1dcb66, 264'h00c5fa3b243e9148e1dcfc27abd9991a2c0c2d25bde9822ce26f344bc9e03f9ee7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{250, 1'b1, 256'hbac4743859e5588409f25335619fe1c7d2000000000056aaa54240b186b1ebc1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00edd7e3fb8581ded7c0961f7365a1a39c6fa301d9728000aeb84c41d918c17dbb, 256'h25cfb4fdade11816359ccfd2001cc2b0e509de9cca0c1aa7eaae719637e11156},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{251, 1'b1, 256'h7eabb2d7d21887903ffba869f353928bd5000000002d3e45954e4b6e21fd30d0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4ca5021a99c50916f997009a2f6addc6cb2a57cada7b1eb72821f66ec353516d, 256'h43d471d4043f8fbb0765c059d1b5386b49a530a626d26d2bed4323c0aea5d24a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{252, 1'b1, 256'h951cd3b90eec711648999d2ca3e8e821b86c00000000574333322ca94097a491, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00eb3a1a9165de050206fa045882f7f3bd06bd02c2e825740d72d8cb2a07f45cfb, 256'h394fa8625004c62cb1c8eea02c3411e6a036b4afe14727d497b31d7251d4a20c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{253, 1'b1, 256'h01ca3636d480cdce6ee63cbe3665c7bd88995f000000003f5d61628138af2b7a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7921badf49f2beba3bc6d696494e7f6c74edc3b722247adbc9cf54d02527ef30, 264'h00a45ef9b623bad9a24433afc7e4e2b25270cf07ab20e29ee822255b6ee8da233d},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{254, 1'b1, 256'he64458ff971279b567c8eb016ac86c39f963cbaa0000000056fbecb71ef3fd7b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3e2c342f84cb36f986b72bd19867c359ad195046ef30ca7549df842d33a51ccb, 256'h5b8bfcfc785ff44ccc2651b893b5dfbc12739cc3973988dbb209cd60f4c1b4e2},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{255, 1'b1, 256'hb15bafa66eaa8c73cedfc9568ac5a41a5b0a45e38e00000000f88ffd117bf4eb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00919eb36b4949e319427b2113927fd40f767c11d2c6a991c558438790959c0071, 264'h009e4bfd8bcca87632071bdc109cd47e45c90f7cbbff3ff05a1591585b2f0f6537},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{256, 1'b1, 256'ha0daa5e1d6fb10cf91937045a9adcd668e53d8d302a8000000000223f8bb456a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e36e3c1918e378f12ccaefe24954c4fb77d8a227f7a234a045c2fa69ec0184c4, 256'h65f7b5def112fd96d3c3ddf3aa5bce418ae5cb7322387b18b5b15e2caa78f209},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{257, 1'b1, 256'h4b28f92a09aff0587c6eb0a61588a5f2d6b1e85955436500000000ecacd385fa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0089674f75b7440869f9de0cdde21ef47003309be9f0ff7f858c6f43a3b9067096, 264'h00d37781ff993210da5470ba8ce3c16a088e58e79d7fd0f5e2d2336443d9b1aeb8},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{258, 1'b1, 256'h1d29293e1f2113a0eec5780d25200ee18779ad86ca0431390000000088a9c6e0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h584c05af98b487e9a0b5dd5e0154d124aeefa55eb48a274721365e597549ec98, 256'h47b4127c6c09077615a921be38942baa053a88b73884dfadd6a745cc9c6fa096},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{259, 1'b1, 256'h3f466438a18ea4e57a572e3ee501d7919c87bb35179a13bc5a00000000023949, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5f21b554fd91ca9cdd5109a00ab3ecb2d8b5137b4fd05c254c3faaa377b3da06, 256'h5d036a7dbebf9351c88d3bbe03991690cb7b67d3b5ca4266eb25029e3a1f75e6},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{260, 1'b1, 256'haa2ef39293ec474361e7562735439b835b55d17b130df2421eb200000000fc40, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6a309780826539059b3b2c9d4315bbb83b4c3afc218d440acf2d01ec0a5cdf83, 256'h5d3ea569a5ad21db62e4bc0b60251e5f65b01158f2c8821973ee6c47cd15fc34},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{261, 1'b1, 256'h1df7127ff896950a28abfee5f9dd0da5da0f5960cfb1d46fc1617800000000d9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h41d51f04d6fdcc5f5cacf88e50e418ef0067f8d854dc991615003f1e49927a53, 264'h00c6f7c10cad03b89460a9794a171f2e10d84982c462cbf075b06738b3f904cc5c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{262, 1'b1, 256'h69e86af97404788bda6b6925dd727c578ada594a03d4975b545b70a800000000, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00da8e729ac23689e868129854fbbde5c9130ebad0e555047f6c4ffccdb0d75fde, 264'h00b693c1a3ccd93e2989f84e77e0ea5983b758f4c1a2a8c4b6219b6b006e9ba1e5},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{263, 1'b1, 256'hfffffffffbda4755bba6de00c2701a0c6fd32c7e4aa1d876140f979cc80f34c6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0793b70b17c7db1ee4f84a0fcc27115355bca4036e33830bddb58aaaf21db1e9, 264'h00b884dc3329f826a3cc1766ab7f67cd31ad17b4d48e81b8641d6cf70400c80649},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{264, 1'b1, 256'h22ffffffffacfab2fac775cbddf678eac83d9fa2dcaa8379ca3af3fb8dd614df, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3ee201732af7f4fb862991d162a11f79fae57233ff964782db1b35b2dee67f60, 256'h78e00f30babf2d483c9e9729c50ac07df9abe878ff8edd3cd7ea3cecc30b724e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{265, 1'b1, 256'ha92dffffffff4bf463c8eca0c62afb2c35c2a592ad8e8e688aa521a258f47338, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h008f2c4f9daeae645deb8237f2598485a7c3ac3b0e0b945641e4f24f59ffe7845a, 264'h00a7f781e40a73cc4f49159ed982ffb264097c5f34382314ba0128a52c9144fd33},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{266, 1'b1, 256'hd0fab1ffffffffbf5c5a0dc94820af6ed2c80b5411be656e273b963141464e36, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h750dad3a83d3c3621a78dcd92f7da948c6fc68d7f0d9603835b2488515c539ae, 264'h00a0736c57503c76c2342e3f13e55f6dfb6637b1fb6ba5caf00b9e540daa7f70c6},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{267, 1'b1, 256'hdf0ffccdffffffff58bc3fac8197329161b5dea9f0043e8cec2a9a631ea38cea, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b3d14a7f7dd693c7fd62d073cb6bc77504431d8a992cc64af774703a981db0a1, 264'h00ab8a35acce773242850c086013869631e99cf9c5378d39d0fe10ca7b504c0cf9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{268, 1'b1, 256'h4d77a2c899ffffffffb8c2d8566f592706ca04276262ff7cfdba0b2ad6e2a6c4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ff35621d420e7a8343d222f18acb46ae5a5a29320f88e2f0977acfd96d701441, 264'h009fc29bfd8a80a24959bd4494de1b3c0a3366131aefef4fe9d33f1f91d118bb27},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{269, 1'b1, 256'heef9d05b88a0ffffffff18a16611a3f3ac44331426f2bdbd5af203e092e61176, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h051291f27408436b4c56cc8993b3891c5c3a4bf3747041b4d915fdccc1c67a59, 264'h00f8d6971a948332617564b4c9581850f8992752f1afe30370a4d36af72376672f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{270, 1'b1, 256'h7e6d3c190be6c8ffffffff27a4b129531bcb4fad150112ceeeeb8d10098dcfaa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b820f2163d1a902e847c69392da7124bc31f56ecad5f73c3db142c9c8220cc65, 264'h0089c527e55e559aa5efb263860fbac04f1ce556f82bcccb49991bc2c575808aa7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{271, 1'b1, 256'h0edd238c04bee70affffffff0ae88780ec5271030a1847cd73f722925df9dd43, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0180c08e97d4fe407c0eab2eb7d17bae60e8ca9ad459e57cdf48389ed9ed9536, 256'h7d5eaeffffba65afbf1ba9ca9bc0fe1181da76e5e41ade8687799b09e9104597},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{272, 1'b1, 256'h4dd115320049ee2e9dffffffff0de268e472eae1699ca5afb5c838313db94bed, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00985f15f0eecc62112817bc234784d60404804ea7dba48f8c09cc02401c4e13ae, 264'h00c73d1bed7077734492c700ede8e6800e048523ef9bcffb53cc79945805ff711e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{273, 1'b1, 256'h1a1109052e9ab4f5dd2cffffffffb1e4604e058f3040a4af85f1f303bd3830cb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d9a5ae9012bcacfc12fa3db623d2099657d4f321460d0135bc731a70478b79bc, 264'h00a5d882aa5cf390737839443ab059d68282064d3d827bfef52fc176d0de60ed46},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{274, 1'b1, 256'h6162159e82cf80a70b34f2ffffffff193b3c777305a8fc809337cb13014edc7a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f070e1285c47106a1ad23a774756a3d3453a48d245401604ef59a96b9a1910c2, 264'h00b43cf52041613dbf8d3a136a0d0f6bce87cd74262224e620f355ddeced20e5bd},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{275, 1'b1, 256'hb35876d301bf4040fac24355ffffffff7fd82e02fe5885a42240d05fff5fc61b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00963a3ae4b0a7ae86047e47f375c7e42de035f28fb430c408d0d815caebefa344, 264'h00a1edd8c2d39f04f99e05a793b7970dfa76f4b1fc0663d308edee9d3ecd077d66},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{276, 1'b1, 256'hc5ae766a399aa8c082a59a4f62ffffffffab6578abad5454b86f0be4e36bedc8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e6adb9139cf47dae0890006732629c8e095c13df370717a42a8bc6e8936678ef, 264'h00a8df8acc7ee7551cf0409e8c1c2fd0df6e7e9b3827e95727fa492c274e4668fc},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{277, 1'b1, 256'h619548e83b2bf592724b244359f9ffffffff7ed41c49517b65795ef980c30f19, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h07662a36a2bb779a276145e78543c360c7d0a22a1749f69ead2788c75750d248, 256'h7c0a4dba499b27cc249a705ba7bbf512a7484b93f9a83ca9305dd49cde6a302b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{278, 1'b1, 256'h2ca970c6acc18b4ad3b023ba01ac4bffffffff4fa0a25f4f35f9b408dd09517f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h36df003efdbec3bf53a2a45248c1e96e60c9bcf10b4f5dfb220744d2da51fc8e, 264'h00e5f103b3a74fa1d0a78e74d604f31889e6637cff2acbb31a70726e72f392d4ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{279, 1'b1, 256'hbd67ed69ca5085f9326153231b96b177ffffffffffb1a4447142406fbb23dd5c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h712dc3233f462b0a37f020ec559bb1a19d879ae36210c75efcb9c071915116e1, 256'h06a981761249cc1929f5c18d6f2a76eef487bbda0c4470bb098b87b91328083f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{280, 1'b1, 256'hacfb85a5cfe484ca5801b819b3e4159dffffffffe10cb294343a640526d5faf1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h10e373d1cb4c05295b63ce7103817b7c0fd096d7c63f65f56d950a61e455c1cb, 256'h44cb5c8270c069ac408a6c9f31ace9229ab6078a36adc465107f0a3d6ddfea66},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{281, 1'b1, 256'h62c18f3f3271e3341a7d3033529b28a2c3ffffffff4e9cf2e8ef755e0953597f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00cd1274f4c89ab194203ccb5c39e7d0bc364537b84b9dd48d922e43e79e4258c2, 256'h42e1fcf72eb65d76b13128d3065daa31312bf9c110f18b4799dce8eccae52d67},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{282, 1'b1, 256'h2df78ec6d8628aeba725a007584b63636883ffffffff0ca2480cb4e3523b2daa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h516c983fe6567ac700f93028da6affc598dfa95391896c544c8f73c96314a0a0, 264'h00bfa56a1833668acfd14899e8cc160b79c5e92a30055dd7c700484f6bfce42cfd},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{283, 1'b1, 256'h07fc58409c7cb5c7169a63d09e4de5120132b8ffffffff1f95f5e389535720ac, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h52279b3df58e2aa7ddaee1e5de155cb75d4f00ec7db74ae913a6ed33dea896d4, 264'h00ef5823ff9977fa492483bcbfc1d0bd765fd6dfa78cc11e658b4984b543e0e79e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{284, 1'b1, 256'h383dfba6e0aa10f820e15e27374c2eb6996baf43ffffffff66a94ff532236f85, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h01c2a04eef5827e7e04eb51802cc3859af6d84fe35aee4da4bc1b0ee154b7ef3, 264'h00dc57a107da6bb12624313660233cbdcc55ff7147ecb3a328af3e86225c89be53},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{285, 1'b1, 256'hc41a8affa1bbbe99587538b31e0b61f8b56ebe58d7ffffffff45e1ee3efb6c66, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1ce1bb1fc78a38d4af211b5fceebd01126c10ceab1de6401e1df1dc495dbf5b5, 264'h00c9b564a0a5b9675eece3cbe33498634e7943893fe16c61ef894bd4be349a6874},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{286, 1'b1, 256'h26fa9d690a2129917bc3520b913f913f1f081bea9aa3ffffffff0fd642c24a4a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b7ae42b36f060c15c6745ea4d8bd91ae2eafe0e196c52cfac4e16ab74d3048b6, 256'h421bc2dcd0854dd4e69a3e930b2cb646557bd68c800c5a2ca7bbb3ddd32370aa},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{287, 1'b1, 256'hb291bf1a8c66adc9def9a0a96da478aa1d09e06797adcdffffffff8fb0460842, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d51dc206df9cfb7198e22b957c644357542264badf5aede3f7474534da0d5b22, 256'h266d172a6d6775963f9ed4fb59065c8f1948c48a51463fe79bbf1b45df7e57b9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{288, 1'b1, 256'h81d64896fa11ee94e49755c0180cc0478de87bf9969ae759ffffffffb4b7f4f5, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f881b3e21684fbf899f762c8fc7c7423a2ad2c276257c99eae86b66ee39e4ae1, 256'h27207d5ccff773b26bf0d282d884b3c3a6724ba06a1671c9f9be8cbe6e3589e4},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{289, 1'b1, 256'h3b88244a6ae111bc752afc8f997cc9ed1f9d4079a0f644f3d8ffffffffa41c42, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2455ebf62b50f958781792fdc705755923a30c0eb7d515a0988c1a14de62caad, 256'h10bd68c881416205bd95a5f2765d69726e0bce5b2a0ec525aeb1bba7d35d8e4a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{290, 1'b1, 256'hbae669421b6378571d97fee160d401bf8f4698bcfa6788a85be7ffffffff6844, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009119d7949d9e4c55e4c712d257c4ba3ab9d657c7e0aa7840091cb2acfb4fc25a, 256'h42524fd0c4ae8b50644cba34f86c21a42ee045ce7c15b4eb817affc78d20fdb3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{291, 1'b1, 256'h1f52ed3bbbeeaa23026b261a17bc00058f2e37cba29772831b7ed9ffffffff02, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h191e716669d84631a04cc085f03b2f1a4f55810f70bebbaf5ee13d68f2598ffb, 264'h0090f208a9f1c27911b5fb8d867bdf123dd601639c2dfa1f6a61fd2f82cadb1361},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{292, 1'b1, 256'habacfdf5c9518bfcd685890b4e11728fe6bb738a9517baacd701149affffffff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h008cc2cab9f257928181c4d3685d544bec0b88b95cbbdb8ad1b0543b46b2414473, 264'h009d1d158dab8e91c68b372ade107aac5c22f8be64463b0c23340dfc828d7b7df3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{293, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h27504e893fd62d0bfdeaa073106b16e8f8d2726a9762529764cfe8fe8a38460e, 256'h21bb0ddff040b7aff8f08a60d5ae1a59472f394846ae4f58c4be0cc8a2a36501, 136'h014551231950b75fc4402da1722fc9baeb, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=136b(17B), s=264b(33B)
  '{294, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h27504e893fd62d0bfdeaa073106b16e8f8d2726a9762529764cfe8fe8a38460e, 256'h21bb0ddff040b7aff8f08a60d5ae1a59472f394846ae4f58c4be0cc8a2a36501, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2c, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{295, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f131f6dddde59bae7b0090a47bafbb33c157ac6da439324a6681bf67f575f90b, 264'h00eccc2fb2c0be318fda9335bb83488bcafd33be82c38318bcf845fd0e5017c248, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{296, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h1101c496d5f8910a7749efff9dc46f68a7fd02d6975fdf15bf90efb70463cb4e, 264'h00de199e46e67d463aa8c752cac8a342b8fe0e9a5ba9a67416c8865c45e478007e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3e9a7582886089c62fb840cf3b83061cd1cff3ae4341808bb5bdee6191174177},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{297, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6e43a5c63ad0bc8d178a745192671c06500f0dbd757c3f2eae65089aaf0d6489, 264'h0082954ff60c3460a27748445525c6cd30701725e1697891cb7f32feed128a3ae7, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h24238e70b431b1a64efdf9032669939d4b77f249503fc6905feb7540dea3e6d2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{298, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00ef4e8b5732f51a4b2547c6581381ccf750bb6d30a07cb758865414d9a45017fb, 264'h00f10247bcaa4ca73d5c9ad4c8a03a60a7f5cfa07fb57437b5a6f0a9bd381d78a5, 8'h01, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{299, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00a973c15a44d2dcd50558e033d242155a29808b87491576566a83821b650e6f2d, 264'h00fc5ecd5482fa591f578308b09f2e704116a375ba1e2837912bae2972d340414d, 8'h01, 8'h02},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h008cd31f1656b21ec27276a533c35bf51d95490bfec57868a9b94433eda4579d61, 264'h00bb2c8e80c45d949bcaf6f0bbc76bc27c95939945052ad1a11014756556c6f978, 8'h01, 8'h03},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{301, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h008cd31f1656b21ec27276a533c35bf51d95490bfec57868a9b94433eda4579d61, 264'h00bb2c8e80c45d949bcaf6f0bbc76bc27c95939945052ad1a11014756556c6f978, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h03},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{302, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h7f77dbb4e500dc9e405ebd9082afa9d0afb5c519fdce252910fcc9202895661c, 264'h00efce51d16a51700a672db8de2af070391a02da1c6a398b7dda94403a06db03d1, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd04917c8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{303, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h6d4f41c9c4c15f02a199264a51266ed793952a7cea79125dcded805ed7a54c13, 256'h50314fa927966b90b6c4e57cb521666fce4cb81b7e4d3550d729fe6dd6bbe5ab, 16'h0101, 264'h00c58b162c58b162c58b162c58b162c58a1b242973853e16db75c8a1a71da4d39d},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=16b(2B), s=264b(33B)
  '{304, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h3bd4a602119bc50cfd05aa395c3c9f753b383bdd9539d27a1a143033fcfcaaa8, 264'h0092d75438eba5af693196d4b7953184e2d649a0845d11af3c7d39e3b1f5449c19, 56'h2d9b4d347952cc, 264'h00fcbc5103d0da267477d1791461cf2aa44bf9d43198f79507bd8779d69a13108e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=56b(7B), s=264b(33B)
  '{305, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h7c981d6870575725427fc84ce6b5f706af6e8c62b4b5f7f72c3ee2860836996d, 256'h29f07476cbf3f93a34e73f737658070642c66d0e34f5d56c715a26b099078413, 104'h1033e67e37b32b445580bf4efc, 264'h00906f906f906f906f906f906f906f906ed8e426f7b1968c35a204236a579723d2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=104b(13B), s=264b(33B)
  '{306, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d75a78cf296b58aeb52faee6a9348385bcdc61f980da8ad6f28654d86fe516e2, 256'h0ce9952182f5f06cba50db8c65aa6f8cf1a32f2a46599c0a2abb4c1402cef467, 16'h0101, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=16b(2B), s=256b(32B)
  '{307, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h0a35a42fb4057e11e332442d73729cdc684e7e0a7875ec933337e74ab1e17de6, 256'h2152e3a6558865d7f30a950c64e9f2e9d2f06c2703d2a1984a79445d3870a1cf, 104'h062522bbd3ecbe7c39e93e7c26, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=104b(13B), s=256b(32B)
  '{308, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h705e0c3ea1ca443a0105896e7af2b891a08243cca510cb5fffaebdd86ec6fc8c, 256'h25d116fcf912e8246a64d5878436dfc958b59d4662a4b227a006876b5042fa58, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd03640c1, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{309, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e322c7aad4a70024c4f80ea373e7e85f23dcbd11f186d55d5a744cd0f459f6db, 256'h71d54db09ec66eeadbedbacfe2255bb87d0c1a737b3d3b1c7b76ce78d6342d7c, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{310, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e322c7aad4a70024c4f80ea373e7e85f23dcbd11f186d55d5a744cd0f459f6db, 256'h71d54db09ec66eeadbedbacfe2255bb87d0c1a737b3d3b1c7b76ce78d6342d7c, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{311, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h4b242ee4a0a37835c590f6abe1af6668476c9c12c15b8aff776c7e7a8a452319, 264'h00b720cffae6423cf47aa375fe3b84346a83b09e0efa245eb89d99b2585451603d, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{312, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f9532aa189138b5e203f8f3a9acf03affa80794f37b647ac289267e8293ededc, 256'h61ac8ac734bc4c7676bbbf57ead50b4981d9bceee0172e947c22c05f4424c9b2, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{313, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h0f2256392bbc44714d5fd698b611b7140c3031845f14f8660baea5ec830088f5, 264'h00d5650dc0f784bd907f41b13936a2d13d0e05deb103efb069f8a771b527322155, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a1},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{314, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h260b66d47b3a3be44364f1fbdd576b824893ce43c78e474db3c1b25106fb4865, 256'h03620b6068877f8b9018efe98191b24cf667053c09ca94da7bcf854bf6924332, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{315, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h30549bef5174962c5650944bbd7833220338e2e31f27775666f7d124d8ed7783, 264'h00f43ee6599a8458c9d786dd50cc676babf489757ade3e267d87bf2654a34adb20, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 264'h00a8ce483b42fb3461047c96ca00d1ab82c81e3d602cfdab62e059b19562bb03f3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{316, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h22283ca6f055439e8540454f63ff02e2e1141d10e34a54737599fae66266636d, 264'h00c8fef97c98fa1160f829b7c1326a069e0bb442428f1503e8cfbb616cd8118832, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{317, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h068f523d44cbb14a249394861c4f417c19dba72f74e1b123b4cbb89c74541b41, 256'h44cd654d2b5871942e8d181f9e38f3946b3a73755a20e68ba555d56de6e290f4, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 264'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa9d1c9e899ca306ad27fe1945de0242b89},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{318, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h123670ccceb86a9d5fce24f070de8dfab093ee66047b17c1d7cca4734820daed, 256'h76495f92804999f894c0184f72235b2db0a7d8ad077427b346d41f24eb2210a1, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h1d109296e9ac43dfa92bcdbcaa64c6d3fb858a822b6e519d9fd2e45279d3bf1a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{319, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f5ab53b565f170a3a83e61dc8cb5bb3a217398f0880db80c41da746d53399397, 256'h3d113d69a23e02aeb2e335b28b85490ace7df18279e2f4a7bd6f69c656fe6763, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3a8a53a9b98a2111e0c5e758a61f57822ead6ac1b9489d7b1bae29dc1dda7a87},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{320, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d0abcee886b680233390f1e6d5ce27056cbfec35ba9231725849a3714b06e828, 256'h5bb11395652a85301cf5110d75d404a1f449ab2ac4767013fd586a9b58114006, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00ac2416840b83e89e188d94463bd19cdc296fb2f891782dbd736b7241d371e890},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{321, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h0f82392f4912bad8f4fcb151b290003174526a8cb27091d38c2aed163040698c, 264'h00dc34e9542d264ecffcd6339963804d68fc8a7376312b8a590d836e1ce1a9e637, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2ec9288261d8fbcda8ce483b42fb3460c908624c8869161e6b15d76e66ec5dff},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{322, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h3b8497a00342aa0ca81408f40de05e938a151e6207a912bc35a13ab8ce8682d4, 256'h75d9d40f07fa88a7418e10d0f92bd10f646016be181c04af65e9ac1858f8e145, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h009288261d8fbcda8ce483b42fb34610470f37567e692db81ce2caa2fe67594614},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{323, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e95914e5d692f4c30724c50a232d432a09664e1d485ecfc3a8299b7007b990b5, 256'h01a21060c529f3776a1df1b3828157dbcd432e84d3ac229585bc9234341788a8, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h25104c3b1f79b519c907685f668c208f63bfd0162312cffe05c2e76ffe7c4ae7},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{324, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00af3e088449e97df3df478c59536965a18598122efc5bb20d23b9f5e41bc84e8a, 256'h403177e836fa23bb3ba2b8fe6005c8d79e1392dc3b726dca4eca14e88c00fdfd, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h61d8fbcda8ce483b42fb3461047c96c9847a30c583c9b9f495591fa1e037b4fe},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{325, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00acaf208d26995e464ebcc54a683b04985c7be74448927e5c15332852886e6d74, 264'h008b182e2468f86cae75d045dc426383d2da3c7e3ab515580f3ff6523f03ce40dc, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00856739764fc50a930e4201325d77815bcf9b7681ed11213a053e816c5df8e6c6},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{326, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h7821e20d3938bbb48240ff48096e928e404ed91eefa37ea7cb2c8f339347b6ee, 256'h6f7ada5c814f0f06eae9516a7848361cc3ac2eb4450a4455743d363f84f0dd1d, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h512c9e1178d280d8464412f2bdf2dd9a7e8065b7ba9216f700779794c9a849bd},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{327, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h009b0ef17c0bd3dea11be2c3358058a1e10b0283108bf79aaae34355c2329e84a0, 264'h00955f5cf7cb593ee756cf4c9f2f0a488a2993aeba923320bfab98c6f72e079d73, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00c9e4be241bd52c69a2486b6d22291f502f64efab87e244d33cacce68672fd44b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{328, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h4ba97363a7e14ce09480bd3b88491a7a501b5d4871b470498abc9a698c069955, 264'h008ce9e198c1d48ec6650d59c15f9e1fb40dc0adccdea6329613e3a9a4decc80f8, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00b0a10528cded5f2b80520ac549338c3f61bbb6f69877aa1b2fe9129c0ce717f2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{329, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h0bad8d9f015770ed8ac654528717734214fff813809b5eb886f87c46d1bac68f, 264'h00c9134ebed0d79a82321cec4c77d5b91c1c7e3c34f6a69cc10140127421b87b92, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00f177b6b48b29de102b6a1921aacd9c94bcec17a59991776cefe8ec63934c61b4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{330, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00ab53f0d664c621138893fc5ee2b26ad2d686bbbb67eda1ee0dfb9609a3f5777a, 264'h00fcf2d72bbd357bea8a1545fd4f162f3faf43bf74666cf23914c7e3d8dde79e97, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00e2ef6d691653bc2056d43243559b392abf29526483da4e9e1fff7a3a56628227},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{331, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h418698cfe9d564e0e5d04a901c062042d864091573f2820f4592d40027dcfe26, 256'h34909e2b92b3cbc595203553121ca46efdda2c23ca990e1e56137365c5a5b795, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00d467241da17d9a30823e4b650068d5c0c1668d236e2325cf501608111978a29a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{332, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00dc0515e400e3527d2785e4a21d105af4cae862b31e07de117f11c9cd8dc9bc9b, 256'h034eef9d96a56c0e74efa10a9f75e2a44d1337e8008175fbb40fe1c700144601, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h56120b4205c1f44f0c46ca231de8ce6e14b7d97c48bc16deb9b5b920e9b8f448},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{333, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h53ff623b312669b48cc8a120b76a811e48a930548de8476d2c4607a5524ce592, 256'h477ae28b239f626067a1d3dee97d769d37b41b184bae95009e401e443e930ef7, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00d55555555555555555555555555555547c74934474db157d2a8c3f088aced62a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{334, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00d2d5348db9d837537c90e930ce35d4cd90e7d7a3460b1384790b632281b98ce8, 256'h43cc7b9a20c8734ac2c62a7d207105f5b2d85c2418939d35e3886f3893cb21b4, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00c1777c8853938e536213c02464a936000ba1e21c0fc62075d46c624e23b52f31},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{335, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00c5fe4159e0b606879fc2a11088d658030ed7fef2e6711aab04869612fd09c3da, 264'h00ac9dc7e198495afc0f43f4de434b8da233d8492cda28db460e8480aecb0a88f5, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h30bbb794db588363b40679f6c182a50d3ce9679acdd3ffbe36d7813dacbdc818},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{336, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h009a72b785c90a695b8e355f5d8fc151046c360d739136241c7fd1e77a0e8b8545, 264'h00a470b4b9a54d1d42956ac43b9c9f2f0f5489da16130b7ba1da38516c912009bc, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2c37fd995622c4fb7fffffffffffffffc7cee745110cb45ab558ed7c90c15a2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{337, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h0081e427bc8f0509b19a14c16e8883b12641d1d68e070c36ab49d1690e5decd061, 264'h00a993d77e9bc0f2b66edc6cd7ca8e32becf32596405622ea2756006deb3e8ac5f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h7fd995622c4fb7ffffffffffffffffff5d883ffab5b32652ccdcaa290fccb97d},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{338, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h756279b4827c83372130d4feab66a4397ed4463ac9ee1dc8adcaddcfcec59269, 264'h00b6323337d89af4208ad8818b67e26f9b8080316bc43fab53d1b3b7cea5db9947, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00ffb32ac4589f6ffffffffffffffffffebb107ff56b664ca599b954521f9972fa},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{339, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00cf9345e850417aa81b01a941a02c5546950c27830841a435f4f3654927c6926d, 256'h1ec53d04954a47f37915dddb48272fe733322d8250783991709b37d87fa296ef, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5622c4fb7fffffffffffffffffffffff928a8f1c7ac7bec1808b9f61c01ec327},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{340, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f95f625795e6cc17b4c28b1ec643c36a34989084aa6a513812c3aa9bec073031, 256'h2b22ce0eeeee9d45cee863c1b1d05381ac8b2c896a2cb17d3e9070d41d68bbea, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h44104104104104104104104104104103b87853fd3b7d3f8e175125b4382f25ed},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{341, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00c3f0aadef8675dc8832a29b397488d6a4fb54780e5967e8b43449498c16ad4bd, 264'h00cb391b545464668d4d0a80b8e283132448a3c0be0abed304cf0839b5920f3867, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2739ce739ce739ce739ce739ce739ce705560298d1f2f08dc419ac273a5b54d9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{342, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h76b920709a9e5dc54a91bd4772ab2593a76f38841dae2880f547c3bb753ae7c1, 256'h5f01e6779d5e3aba75997bcf7e3f320868ba8f0bc1210ab80b42760a6a701206, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00b777777777777777777777777777777688e6a1fe808a97a348671222ff16b863},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{343, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e3895147f4e36a13c3483ac00c88a78a8ffa42478afc2e9d8386205b0b1df8b2, 264'h00b4156b56ba217b1ca08bd77f819abb52d742f6b2f7d61353e4cc5663da487317, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6492492492492492492492492492492406dd3a19b8d5fb875235963c593bd2d3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{344, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e733999ce348cf7b363dcf931953cf1c247c3a887408c064b9791c178ad35029, 256'h0b0849329da7008e6a2d00142883f8041b9917528fcc4c5bd3f795accff28eb6, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00955555555555555555555555555555547c74934474db157d2a8c3f088aced62c},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{345, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h069b66f716902cbd51dadff61644ac74c6a35e8c776ea22c9c3492d1d3faa2ec, 264'h00e4905cc480bc967ce389b82c8e6692b159d3fe9a268bfc12010993934d7e24dd, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa3e3a49a23a6d8abe95461f8445676b17},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{346, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h009543bfd3a0b678654fc65458e3e62269b30bbd2a40282d92058c3311a61bd885, 256'h333d78221d9aa0a9663a5df5123d95c3ff4a02606278666179e33c94fe1e0cd1, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00bffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364143},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{347, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00a6884e6218642518a211f67b03aef6a84d3b32d18eea445b31913e8a1a00f4c5, 256'h31a318166cfcbce34307572eb823edc5d0334c5e5373af4e832e730047996aca, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h185ddbca6dac41b1da033cfb60c152869e74b3cd66e9ffdf1b6bc09ed65ee40c},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{348, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00bd4c6f9ab363a204fd1abe0f7158b84417cca2e0d355277ddc17cac22abdbc2d, 264'h00c66469bb8e8e04186e81a2b693cc2121ef22cb61803a2b4ebe1a3e0d367b295d, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 264'h00eaafe4ce77ccd9137f39edc5370d26b73f4dc6ceadfb40a488b2dc6c93f1993c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{349, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00bd4c6f9ab363a204fd1abe0f7158b84417cca2e0d355277ddc17cac22abdbc2d, 256'h399b96447171fbe7917e5d496c33dede10dd349e7fc5d4b141e5c1f1c984d2d2, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 264'h00eaafe4ce77ccd9137f39edc5370d26b73f4dc6ceadfb40a488b2dc6c93f1993c},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{350, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e1815bb1653b8146a2e9160fb0e946112b8994b9d90ef8a36a8ef2ba187b705d, 256'h11b344caed87db94b9c9eab8a5e3277a9aa46b31768cee5406c3cbcffce0a945, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0, 256'h33333333333333333333333333333332f222f8faefdb533f265d461c29a47373},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{351, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2be9265c148fc61379ca147e651e7f0a1c602cdd66f70b4b6ada2e83f56c1a71, 264'h00f5e1ede0139baa93af588cc7ec1b479b91d230c811575cb143af12c631d16a61, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{352, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00af3b3f73a409ffa51b10f3cdfa272d9b42358ca9aed2840bfaf5bd67e61fd1c4, 264'h009d07371ca919a069e46c473e6e45b2f2cd019fa21f84d0abfa285be5513781fb, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 264'h00b6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{353, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00e155240c3be314924ed787354325fdc3dcfe46d603798f2491152448e0e413b6, 264'h00ce1124313eb0048292f6edf9f248ff9624936e41be6c93dce2df9ab7997289fc, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 264'h0099999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{354, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h0087d4de4ed890da42d7e11a95e56070c95901500c53dd55b62952679884d2598d, 264'h00df8a37ce6d8f86f4e8b3580d6e6a448520cb740888a3b0eac92bc9a2f1589b4e, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{355, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h008c03d72664214f3bdaa6a2e1003b14864000e5993b41b71b68cdebc4a08f628a, 256'h4a490efc9172983bec203e6096dd9778bec26f6e443e1dde67060dac18ca2440, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{356, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h1ae8bf7b21b3ae00fd01d19b4f72ae6b47bf752edf476cc5cdfa1c2345588e71, 256'h54dc306165f4f907802478ed2aed41ec54ddf870bc62c2c373971194308411f0, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{357, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00c5dad21249273cd72ad06943b4e3be0822595bf9fa0459223d27354dea24179b, 264'h0097340abb326afd1eb6de5e525a23aad4929f8a09244c972841a0cb76680ff060, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{358, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00f2c6643bf373a0812f993cd616993551d7bc7826d3d6bed0918ed4998b74e837, 264'h00d7160a452dd2c8d3e5f4f80a1efbc33793c35d6e243e9dfe9a39e26dfb7a1b9f, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{359, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h3a1bd608d3187c684d8d461a5406e2b86b09eedc5d2dd28fcc341bd2d483a6d8, 256'h5e3ab9d9e79ecb7e43135782ae60b12ff69b3349c1819b4ab27b738c7f803595, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h0099999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{360, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00aee2e5aa96d31bde8b0ec1e71d79e721c5fb094eba49d61dfba6e636a77b215a, 264'h00af3534fa210143ce3cecc5bfe1e0b136ab6811d662376637efe1eddd212b6ff0, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{361, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h00db0dc63f6dfff9b2564498a2423449cc5d894222ddda86eabd6d2bb2549d28d7, 256'h5b5bc20153ef6a2649dc6f116e6ca5c916740a9a645618003a5a448eee928fcc, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{362, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 264'h0082a004a2ff4aa7c2fd4c71bc88a4ee16d75c11f5ad8599a6eb41ea73e49f80bc, 264'h00f360abc795b4b21b46584a1bebc41720df51a25044880f287c5e5d83f83c1d20, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{363, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{364, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 264'h00a8ce483b42fb3461047c96ca00d1ab82c81e3d602cfdab62e059b19562bb03f3, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{365, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{366, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 264'h00a8ce483b42fb3461047c96ca00d1ab82c81e3d602cfdab62e059b19562bb03f3, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{367, 1'b1, 256'ha7ffc6f8bf1ed76651c14756a061d662f580ff4de43b49fa82d80a4b80f8434a, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 264'h00fc0f737a79d525eefe3c940c162173cc6fd9a6d5cc5017754026c4113d0f15cc, 264'h00894d6fb59cc79199b89cf12b556ba49f8623b66da8c11a55e267e3318497688c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{368, 1'b1, 256'h5a7a8ec92299354caa012069a923d56d0043b22408fb36ff8cd0ecba3aacb0a4, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h76bae33ffa376b496bde93c7748d50a3a8b73bac045e54c40c7fcd344a10fa83, 248'h3e25a20716a902d524d656ead090b7bbe1ac25ff71269d7038d4b08db5b1d7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=248b(31B)
  '{369, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h016e2dfac600c8c994c0bb815b1072bb5bb680774121d342f93fe0a994f72c09, 264'h00c378944de05aaca70c71ed9a7fe4eed2b36ab3ddb4b32d09d53eebd91f2f9217},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{370, 1'b1, 256'hf3683c9e3da9a7f90397767215345efe3be07565f14ab80d102f50644b98fbfa, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 264'h00a33c4acb033f3d0d50d244249a1277448b6a52f524e30f4b73d595fb955e9247, 256'h7f31b50c698a971c8fab98521ef3a1d6fa483a676230467c8af3018452bf1de1},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{371, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h091bc829be861c20c4bb877f0da205b3911584708ddeef580ae46691b245b99d, 264'h00c03bb5e77a8fad94736775f31ae381015a93973954b2f3e541457fcb05bccb5f},  // lens: hash=256b(32B), x=256b(32B), y=232b(29B), r=256b(32B), s=264b(33B)
  '{372, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 264'h00fd6a7eec40d1062b9a4a7af4817b3ea8cd21596d6dc228b287a21b647caab29f, 264'h00ab861672dfe3b428c26e08f2f7ca464ad3e966bbf62931408ed1ce2735bab62b},  // lens: hash=256b(32B), x=256b(32B), y=232b(29B), r=264b(33B), s=264b(33B)
  '{373, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h53ebb6debd028f195c039ef4e04276adfa2d9551a6e02d2c4143907ec889e6d0, 264'h00fa01a27240dd63aff235cd9778c90a7c25c993791cda584fdcca1a979f5faf54},  // lens: hash=256b(32B), x=256b(32B), y=232b(29B), r=256b(32B), s=264b(33B)
  '{374, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h60ec4f23f1b2c0b5acae075bbf09be76ffc978aa4d354d309746047a69c43ddd, 256'h798c3df3ada3c91845272b9573e70e683d4e49d90a51f6ad047e24da19355d3b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{375, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h4457c32fe6bf74ee82ff8a38b8076b48323769f3b7970f419352283984dde081, 264'h00c6380b3ed90ddba62394c19e02a3b8690d1615dd1120c0fe67b86e7961b8e7d5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{376, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h24820a985bc72c8817ffdec275db7406ed5b897fff0b713d98a721a42bb4c6d4, 264'h0094f1397d1e577fd47cfed7ac01f2aead6888863a3f8ff21f00c34c41e840af99},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{377, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h1ed4e5132e4b11268ad55b9a4b7a54ad3e028976bbe85fef2e8cd0a3e4362c70, 256'h1d1ce94fd8ffda6df3c307150a98719f276381b0c9d261fba7feba37b402394b},  // lens: hash=256b(32B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{378, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h4f030196e9a558b5af5557c7347d132b1308b3a1ce88a6bc6bf566ed22b5da78, 256'h392ddc6e83f995a0030856ecd0822449d8dac2bead6d269ef4b307d535dce238},  // lens: hash=256b(32B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{379, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 264'h009eaa256762ee3d5d3ed269a2907c4a836c92073918be335469e25743ea9ba0e1, 256'h2c70e1dbee671e9bbd6b68695ae40d58d11ce82592cf9824914a1d8d9e429fcc},  // lens: hash=256b(32B), x=232b(29B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{380, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 264'h00db965e2d0d25c84c30ae8a3e31f12b55b8784b90f91d443a70f2c7cb4828f5bf, 264'h00aabb284a7715095cb11714ec76779c08ad5496d8870e2109467a21093f0b8bca},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{381, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'h58675835add3dd65f25c76b02545176c37a840748fb64a16b8bb113e361cf55d, 256'h3b1e25552a5c35732f33735f4dc6f50f947bbecb734599a987f1ffbf86b2842d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{382, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'h786a687776da9c185afa16f90a596f5ddce3c2d3caece0344101be24581b86e1, 256'h75b13da23be046d551c68b54e72a990288dd73099800705e1a854366662b950e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{383, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 264'h00cfce7188667568bd7d5269a75bef42aa360705db5232d189adcf2323036852bb, 256'h5d06871c28d89198870f94264ae11744d254682e06f154332f976b803da8a1a2},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{384, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 264'h00b21cc81843c74779fc5ba9fe1b0d5e7173f696c6e91398cf83a31bc735b6050b, 264'h008945e8711789093c80fe6cec3947cc9c36ffe2505f1ef721bb507e05c9c07bd2},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{385, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 264'h00fbc5087d1e6bbc32dae22a837d03151028ac69ad71e66e5fc841de0548c06dce, 264'h00e2dfa5e56de28d72d0e770e7666033c42431bcae1fc6cffd9593d54cbcfcfa7c},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{386, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h5ea780b73ce027c03ff81e1b26e61076c8944a835d349cd757ece0c4ddf1da24, 264'h00bd9b87db26158d5b9132bb0f3df54a2ab6c9ae9a4e0b8496a539ab4ab588ccba},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{387, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h4618f1a11cf8cbc1966416785c3149f75a71ae256d445deb31008d51ba6088c2, 256'h408087725dd6ce18bfb7493a5460b54022245e5dbd731ed6d35db88a51d2ba6e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{388, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 264'h009d9cdb94e5e9a66bf8eedfdf9f1af43713bb05d880dec89aec21631958970de6, 256'h732932649bea35f11dfe0926618e4f091c1b264ca128a9eef14e6d94d7c9f207}  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
};
`endif
