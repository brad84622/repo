`ifndef WYCHERPROOF_SECP160R2_SHA256_SV
`define WYCHERPROOF_SECP160R2_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp160r2_sha256;

localparam int TEST_VECTORS_SECP160R2_SHA256_NUM = 66;

ecdsa_vector_secp160r2_sha256 test_vectors_secp160r2_sha256 [] = '{
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{116, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=0b(0B), s=160b(20B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=0b(0B)
  '{120, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h08f8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h35a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f93150, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c376ad},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 152'h0af8cf160e6cdee66be28cc2e341d85210f931, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=152b(19B), s=160b(20B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 152'hf8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=152b(19B), s=160b(20B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 152'h37a47217e8565667530eff75cec5615107c376},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=152b(19B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 152'ha47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=152b(19B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=8b(1B)
  '{138, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'hf50730e9f1932119941d733d1cbe27adef06ce30, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'hc85b8de817a9a998acf1008a313a9eaef83c89d3},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{153, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{163, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{243, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h39b0c99df627abb063501b93bc0ec2f9fe1abac9, 160'h01e957fe1c54b5ba221f79b64fc2763fffa80524},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{244, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h2ab314be8a53a6af98e60e9378ad5194a6306629, 160'h60101c49dbbcf678851f678562bb99b0e983d011},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{248, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h53f4103b4ff5f2b04e60409b712b24e52d446bee, 160'h5a0a9c4e5ed87323e7a2f8964cdd05aaca8623f5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{249, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h623a961ae133e8fcc433d41afbc7d479bbacf5a7, 160'h120f4662c44fd860a09057d016ea22f59c9ea48a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{255, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h55a270df082a4d6183a4b6ff10a737e02c48b4b8, 160'h5026129206b77d6b0de92147deb0d0ae7c2260fd},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{256, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h6d84f406773166c41bb442f5af04ab9858df5604, 160'h6aa89196cf9bfe8dbcda618438dc717c8fdc0bc0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{261, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h25952151a5fbe15c4184a0b1f212a8710f51d665, 160'h63c69705d2e525b5533bb545550d421f65a811fb},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{265, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h5f1614bd3ed8ff1755186b3a16d0b46c98d4363a, 160'h70fed0fc130a3e15086d3dd5150b452cc9234dc2},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{266, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h7579791e611efa8183708f49f474db39e729201a, 160'h671ead3c5c8a57b90ce81cafea1cc7ac5c60018c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{269, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0ecdf9992b5ebbee6770dad3aeefaceabc6106ee, 160'h5e849ff0607952682b51c8889d4b1dc0371f47fe},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{270, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h178bd60ae5c02fe00f058e4174535e62caf9ab3d, 160'h631242e73ef54d6e44a5adb7a1119e0467b52e50},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{271, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h755e6da6c7aebfec7169771d70aba265bbbd94b7, 160'h00c19262b7cb5e3be6a4128e54b8ef756f3c9085},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{272, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h7ec65c17c976fdab34e41858e39a48da52168e87, 160'h39df46e7912443837e38dbd210679ffc2be55d99},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{275, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h46591cc99953bc95bd791df1d49852ff4d155933, 160'h719ff20f870dc699c20be7add0701c6ef9f47c28},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{278, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h42c1dbc859090702b337f06304c32855aa032d58, 160'h54eb0ee6de7a6a75dbb3162a320d02433706fe5a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{280, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h6e4fbcfa8f008eaef72bf80224575cf6e0d5a6c3, 160'h1ebe3f075dee784663ec14b687aa54384078b8ae},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{282, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h72526c3ead0bcdf74e527c5498cf1b1df7d8524e, 160'h0b297ed48051140ca2ae592da02dd03e5f25ad84},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{285, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h758a02aa0f79ff94b7b56086f803688072aa25a8, 160'h281a5a69e4571646333cedb80ed565d11a30f964},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{286, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h2660d3799b942b3e300bf7197f79724ddcb1ce47, 160'h3759b27452ff2465a0a947a904d3812e31405362},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00fa19aff61dccb4982a520c4a844210d88245e643, 168'h00cad5c9f87432f65dc9609b50ae80da751a86bd32, 80'h351ee786a819f3a1f4f5, 80'h351ee786a819f3a1f4f4},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=80b(10B), s=80b(10B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h0dd2d6ce794df00949356bda4ce5933b41ebe45b, 160'h71a799413369c351373f18f66ee5ec3f08986c91, 40'h010000538b, 160'h46b6470dc8b43a7f5fe139ec959eafa683f28f2e},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h74151122fd301dec9139e1277de1063810fcf9c6, 168'h00f1797e4233303f7279e8bff017466a2963da7b53, 8'h03, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00af1ee8e681b5db8479ad6d2c3cce1bb6da8c87c3, 160'h427c7f8dc4de05c78a0ffcf5412ef343bb137e12, 8'h03, 8'h03},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{302, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00bebde6a1518a38bcb7fecfb6e70d92ec5de9e2fc, 168'h00931816f21cd2ff7c7317aeccf50a994a6fb44c71, 8'h03, 8'h04},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c7a2767e0ee2fcfcfb9f5956728977d6cb976a37, 160'h11627527eede9dad36f80302c1d39e5707674107, 16'h0100, 160'h4e9d3a74e9d3a74e9d3a8539de479664630141b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=16b(2B), s=160b(20B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h32c14d92c5bbf6e3440c4428bece01c77c4c847c, 160'h3cf05f2e5c56e67c8e583d982b6b4ef498c1cfdb, 56'h2d9b4d347952cc, 160'h6b725fdd61cad3a932f93b73e8fb939d7b7f98a0},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=56b(7B), s=160b(20B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a9309d2aa0520e82039cac944ec6ecdf2f830889, 160'h4291efe0efaf29d95e041b1a423a3b4f4d30c507, 16'h0100, 160'h3cc5990d6ad0679254b205b6210dc1204c382e92},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=16b(2B), s=160b(20B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d500ef5c55e6df67dcd941dad4e138ecb5ff7455, 160'h7d239fc8d9d3da2b799ed6c51f2f542f650eaecc, 104'h062522bbd3ecbe7c39e93e7c24, 160'h3cc5990d6ad0679254b205b6210dc1204c382e92},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=104b(13B), s=160b(20B)
  '{311, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2805fbf5352896e2fa4d0ce04a1e46a1e0a54958, 160'h7d14fdd85792bce2592ec6e3adfab1232a1e1eeb, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2805fbf5352896e2fa4d0ce04a1e46a1e0a54958, 160'h7d14fdd85792bce2592ec6e3adfab1232a1e1eeb, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h300cc0a40c609362f3f20b7c8e57a8f99e592436, 168'h0092a393c1bd3cd2792ca45b8bd56e4f7186817a54, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{346, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b126e61fb24c9932a12c50a14844887677276bca, 168'h00d4710b84ef34a8b28e290179e864ab350c761785, 8'h01, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{348, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e0c8238a5ab89f192a0190821b958986103d0966, 168'h00bd64baf7e2417212d99b4a899264e122db67e99b, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 160'h333333333333333333333dd2fb1aee6b63ed2048},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00ad4577f7f3008aa5ebbe149509ad3de4b7bac270, 168'h009f1a6ba48149bde27ebf3a8fab4b8483676b4c95, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h008779d9d40470df9c4b6c53c27330a0f0c748c01f, 168'h00abe5c16182899fe3d702ee89bb14a51aa8ff6cc7, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h666666666666666666667ba5f635dcd6c7da4091},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a7afd930bd9f9392483245ccd628be428e0f6555, 160'h36c945fee505c5fe855187ee725402995cb0e701, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h6db6db6db6db6db6db6dcd9f87cbfee61f45452e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h45fb936471ddf35059c571f794b7fd6f23f752ff, 160'h3fa9603f8c5a370da68f3f812802f0da5d21af74, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h0eb0f1bc9eaf6ad85b2d94e5e1b53937df61a288},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h49d0064ca551c15fac3f13f9cc44a8309c31e721, 160'h3d403f3bee9ceaa243e492cb9a8f83e92c3c11b6, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h491a910b75f57a4cfc2fa7c878c0a23a725952d5, 168'h00aeeb19e0aba884da4cd64574e785ab9323d0f681, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h666666666666666666667ba5f635dcd6c7da4091},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0099704a8b543c9ee06a913b9476d6e1b741e28368, 168'h00df8cb71743ef9903231dcfeadcacb4e640192397, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h6db6db6db6db6db6db6dcd9f87cbfee61f45452e},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3a81a3afa818e6511baed5c8d52c617223cd3608, 168'h00f3f13a8c30bff4cbfbad5d0789f8e12bce995b43, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h0eb0f1bc9eaf6ad85b2d94e5e1b53937df61a288},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{366, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 160'h46f1a7493b131f3c6032e9612b8e1bd3d1a3104c, 168'h00e3cef3c8020c277ba45bc93a9a364f07eba8302c, 160'h6d8624bff7719b53dab811bdc0e434a5e9f02e8d, 160'h0b50e6dce0f5c1a757290eed8df0aa8092b2ff90}  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
};
`endif // WYCHERPROOF_SECP160R2_SHA256_SV
