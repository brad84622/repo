`ifdef WYCHERPROOF_SECP256R1_SHA512_SV
`define WYCHERPROOF_SECP256R1_SHA512_SV
typedef struct packed {
  int           tc_id;
  logic         valid;  // 1: expected pass; 0: expected fail (zero/oversized)
  logic [511:0]  hash;
  logic [255:0] x;
  logic [255:0] y;
  logic [255:0] r;
  logic [255:0] s;
} ecdsa_vector_secp256r1_sha512;

ecdsa_vector_secp256r1_sha512 test_vectors_secp256r1_sha512 [] = '{
  '{1, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h5f85a63a5be977ad714cea16b10035f07cadf7513ae8cca86f35b7692aafd69f},
  '{2, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{3, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{93, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hf1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c00000, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=34 s_len=32
  '{94, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb20000},  // OUT_OF_RANGE r_len=32 s_len=34
  '{98, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hf1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c00500, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=34 s_len=32
  '{99, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb20500},  // OUT_OF_RANGE r_len=32 s_len=34
  '{114, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // r=0
  '{115, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{118, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2678f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{119, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=32 s_len=33
  '{120, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f98140, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{121, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34e32},
  '{122, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h002478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{123, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0078f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{124, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h00a07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34e},
  '{125, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=33 s_len=32
  '{126, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=32 s_len=34
  '{129, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // r=0
  '{130, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{131, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1cf49f6d858ac900a7af177222661ac95e206d32ee63020beee955ca711, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=33 s_len=32
  '{132, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d149f6d856ac900a7af1772226e7dea086b8a3f1dc48ad29689c965c6f, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=33 s_len=32
  '{133, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdb870e2fb60927a8536ff5850e88ddd95b3a64cba0446f9ec3990bd467067e40, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{134, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdb870e2eb60927a9536ff5850e88ddd918215f79475c0e23b752d6976369a391, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{135, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdb870e30b60927a7536ff5850e88ddd99e536a1df92cd119cfdf41116aa358ef, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=33 s_len=32
  '{136, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=33 s_len=32
  '{137, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdb870e2fb60927a8536ff5850e88ddd95b3a64cba0446f9ec3990bd467067e40, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},
  '{138, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c3a41688548eb315e94effca0efd1ffe0a13467061783dde1cce167403},  // OUT_OF_RANGE r_len=32 s_len=33
  '{139, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c5a41688528eb315e94effca0f835208aec517335790ca4896d5502961},
  '{140, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h5f85a63b5be977ac714cea16b10035f0bfc6fca393d12e237b7beca62e4cb14e},  // OUT_OF_RANGE r_len=32 s_len=33
  '{141, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h5f85a63c5be977ab714cea16b10035f102e001f5ecb98f9e87c221e331e98bfd},  // OUT_OF_RANGE r_len=32 s_len=33
  '{142, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'ha07a59c4a41688538eb315e94effca0f4039035c6c2ed1dc84841359d1b34eb2},  // OUT_OF_RANGE r_len=32 s_len=33
  '{143, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2478f1d049f6d857ac900a7af1772226a4c59b345fbb90613c66f42b98f981c0, 256'h5f85a63b5be977ac714cea16b10035f0bfc6fca393d12e237b7beca62e4cb14e},
  '{144, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // r=0, s=0
  '{145, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // r=0
  '{146, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h00000000000000000000000000000000000000000000000000000000000000ff},  // r=0
  '{147, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // r=0
  '{148, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // r=0
  '{149, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // r=0
  '{150, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // r=0
  '{151, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hffffffff00000001000000000000000000000001000000000000000000000000},  // r=0
  '{154, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{155, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{156, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h00000000000000000000000000000000000000000000000000000000000000ff},
  '{157, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},
  '{158, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},
  '{159, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},
  '{160, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},
  '{161, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hffffffff00000001000000000000000000000001000000000000000000000000},
  '{164, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{165, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{166, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'h00000000000000000000000000000000000000000000000000000000000000ff},
  '{167, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},
  '{168, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},
  '{169, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},
  '{170, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},
  '{171, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00000000000000000000000000000000000000000000000000000000000000ff, 256'hffffffff00000001000000000000000000000001000000000000000000000000},
  '{174, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{175, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{176, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'h00000000000000000000000000000000000000000000000000000000000000ff},
  '{177, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},
  '{178, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},
  '{179, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},
  '{180, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},
  '{181, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 256'hffffffff00000001000000000000000000000001000000000000000000000000},
  '{184, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{185, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{186, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'h00000000000000000000000000000000000000000000000000000000000000ff},
  '{187, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},
  '{188, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},
  '{189, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},
  '{190, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},
  '{191, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 256'hffffffff00000001000000000000000000000001000000000000000000000000},
  '{194, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{195, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{196, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'h00000000000000000000000000000000000000000000000000000000000000ff},
  '{197, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},
  '{198, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},
  '{199, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},
  '{200, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},
  '{201, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 256'hffffffff00000001000000000000000000000001000000000000000000000000},
  '{204, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{205, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{206, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'h00000000000000000000000000000000000000000000000000000000000000ff},
  '{207, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},
  '{208, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},
  '{209, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},
  '{210, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},
  '{211, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 256'hffffffff00000001000000000000000000000001000000000000000000000000},
  '{214, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{215, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{216, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'h00000000000000000000000000000000000000000000000000000000000000ff},
  '{217, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},
  '{218, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},
  '{219, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},
  '{220, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000001000000000000000000000000ffffffffffffffffffffffff},
  '{221, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hffffffff00000001000000000000000000000001000000000000000000000000, 256'hffffffff00000001000000000000000000000001000000000000000000000000},
  '{230, 1'b1, 512'h5f254161af29b81dd51085800b0d053e358ec7006384d8107627aa4bf841bf84e0c85418a7976a1088231175d964c161aaf90e63ca0ba7e9d455b8e80c77bec2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h64a1aab5000d0e804f3e2fc02bdee9be8ff312334e2ba16d11547c97711c898e, 256'h3c623e7f7598376825fa8bc09e727c75794cbb4ee8716ae15c31cd1cbe9ca3ee},
  '{231, 1'b1, 512'h0000000001b99889c891f2468c618149cb6865b933cca31eddb353de09746b540616ba69c5f5ff992c6d6177427daf1cb46a4c5c08625263a615fbf3eeaae178, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3a4f61f7f8c4546e3580f7848411786fee1229a07a6ecf5fb84870869188215d, 256'h18c5ce44354e2274eadb8fea319f8d6f60944532dbaae86bfd8105f253041bcb},
  '{232, 1'b1, 512'h7800000000c52e48c315d5276f18d994c345b5805aa02872c29105d1bf75f152042a782853b4a3850822714434fefe3db00a19bc7eb84029869a7c1dca47ce71, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3fa9975fb2b08b7b6e33f3843099da3f43f1dcfe9b171a60cafd5489ca9c5328, 256'h985a86825a0cc728f5d9dac2a513b49127a06100f0fc4b8b1f200903e0df9ed2},
  '{233, 1'b1, 512'had9a00000000987c9531c475b0236659fdd3dd795473bafb8f0753bcaa4bea4e6418f79cba317764c48fdfd9461986dcf668f250be9ed2b7b75afaac70ccf0ec, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4d66e7ee5edd02ab96db25954050079ef8de1d0f02f34d4d75112eaf3f731240, 256'h6292d1563140013c589be40e599862bdd6bda2103809928928a119b43851a2ce},
  '{234, 1'b1, 512'hb3284200000000930b8b98132341f68419e3262a7f2b8d60cfee7e1e364b36ed4f000bd5fcde187cde7397820b85a174025e4d54d70cbaa80d160fc9cc72d56d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'ha9228305f7b486f568eb65d44e49ba007e3f14b8f23c689c952e4ced1e6cf91e, 256'hb73c74d28bd1268002bed784a6b06c40a90ee5938ea6d08f272d027e0f96a72c},
  '{235, 1'b1, 512'h3bf2ef06000000009638300311c31a5caa29197ef0d079767e66e50824e8d41e5a36f593539a6c0ce102a92493c18061c70eefb94903831d9b8ed3291d1b9829, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3fa39842bfab6c38afa7963c60beb09484d4579fc75ef09efff44e91bc62ca83, 256'h5612add1924f0285ace5b158828e2b32ab2b6e7f10ee68dca1cc54591fee1fec},
  '{236, 1'b1, 512'hef200f1a5400000000399e032faaf4b3c32d804555abf20471a3a18dc46f3917eb9072220b5d5f994d27b221346631c47eb579d69cc5e438b7e7b963bca9d84f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h06c04b02edfeecd8620f035ea4f449bd924593e86e5288a6f22d1923b0e2e8a9, 256'hf666718e6fefb515bb9339d29cc0e58cfba89d605ca0066bca87f6a3f08ebcfa},
  '{237, 1'b1, 512'h7f12580858d000000000055d6877381f726e0a9237d1c012c9840b5b3fbeb6f43027bba37a94ba5fc0dbab436b88d4a7cde6aac151b06214a00cd8fe5f0bdef8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1ddd953c32a5f84109cd4d9ec8c364dd318376ff5d228211a367483077d63880, 256'h563dba4845de762baf04910618d587e0dd0c97dd1c9785c24ffdf2f8a660abf2},
  '{238, 1'b1, 512'h6b4185d1e7382000000000c86f684e5386df6f2e7e1dab4d1be30ccac1ea33d4e82d455b12857120cfb411b75c8df08758216dcb774dedf1438bd137f831b27d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h9fe4ec4831ef4945f100d5d35a2e6312411ca5df6c900ca60690f2985d553482, 256'hc674ad5e1bead2f767c9248e444452a4a8530dd47246cbbc968da865bdf212b6},
  '{239, 1'b1, 512'hd40c1a66696b7a6500000000ebb22b0b1f80b394770ad61c5c42ff0584ed4c84a3d185d3c07725f0d3080b451dad86945cc9b0801c01e0b6b8739ff8ec36df22, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'he8703d6b16a79fc2ab3653cece29d06f65dd6f2c230cb08ee30c5517407d75db, 256'h8cfeb87b8e95ddacd638b37d315393c5005f3ab8bba0cc1cd1a050829b775bfb},
  '{240, 1'b1, 512'h68481d736990000f3d000000001bc2164f3bf7a43f3c7f23a875b84fcc1d1395c9bc3eec02e9aa7d38f4462d5734ca53f0db4e46498d1b8c9f9f4c92f4fc0532, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdef608caf1f277d71403009f209c1d7eef11aaa7920397fbf429b8146181aece, 256'hf3b8f2aa5b3df9a8b37313ea66ad5b74673f3e8614ff471b1eb6773217511fb0},
  '{241, 1'b1, 512'hcf9bb31b573fa12e7e51000000004b37d8761e5d50f214b30bc2b134bc7e0e30653b8debc737a21392357313d13e08eecfdefd8d37bec92b680a84f5430fb57c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4f5d08e8d936ce831d02d6b23fb8fce0e0750101af3ab9c3b28636b95a5e24ad, 256'h6f034480553bcecac221f8be8288163c55492e2e56a88f4d0341b61436a0a6c0},
  '{242, 1'b1, 512'ha678a93e12f88e59d6307e00000000bcef462484d98a07578e5106f6b5e6cd1618aa82e3797b4bf519cdc4704616039255cb3f05fc8b93e4a48e2c4cd5333450, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hbdd822bfe3733d9f4b88764fe091db2e8f8af366e4c44d876bf82e62bd48c7ee, 256'h7fbf7750c5dc849a2c55dbdd067806f869652a7b3a57baa4733781d3128f02de},
  '{243, 1'b1, 512'haed2cc5334773206d7170bca0000000081dafcdf0acf2107d7c016b54b1c0ef3663c5ba78277a328ae547ffdf6ef2e385a374d9355022f24dd05ff9b357e5039, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1c4fc02961b7f4245566b410bf08f447502ea4f75b15690344681efa2edf7b4b, 256'h7d63eef119dc88bc4a1b2c43ac21cd53892443661f8c3a97d558bf888c29f769},
  '{244, 1'b1, 512'hfeac570e6cd1481ff79f34cccc00000000eb127fae412cf598abaa6550b4f5f2e1537dd5c5d6c57b0b52c103ec0340c9e292d0a263d74e44301efe65d505ff9d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6406f2d249ab1264e175476ca3300efd049fcad569dff40b922082b41cc7b7ce, 256'h461872b803383f785077714a9566c4d652e87b2cad90dd4f4cc84bc55004c530},
  '{245, 1'b1, 512'hbacfc820b1f513e6a157534762b6000000008ba56a4c814c4c12a828e658c8f7d0453900871cece52dca13f4f1df23685d1bd43488e2acdda903b2e0f72b9d64, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h415c924b9ba1902b340058117d90623602d48b8280583fb231dc93823b83a153, 256'hf18be8cdc2063a26ab030504d3397dc6e9c6b6c56f4e3a59832c0e4643c0263c},
  '{246, 1'b1, 512'hf9f58ffc6e2662f4992e06774f928d0000000084b7ca7f7b6fb750919f466be3366746484849f67645a424ce6009fc560031052d0775f47984d3a4727776b916, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hd12e96c7d2f177b7cf6d8a1ede060a2b174dc993d43f5fe60f75604824b64fef, 256'h0c97d87035fcca0a5f47fe6461bb30cbaf05b37e4211ec3fcd51fc71a12239ca},
  '{247, 1'b1, 512'h5f6f67fd931001c593ff6f8e5ea8faac00000000ecb4ce9ec81a128cb55bba07a9b186b28f7e787f7bfb7ea32d9047b830a99f2ac4144ee3f6e07ddf00e68646, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7df72a64c7e982c88f83b3a22802690098147e0e42ef4371ef069910858c0646, 256'hadbaa7b10c6a3f995ed5f83d7bda4ba626b355f34a72bf92ff788300b70e72d0},
  '{248, 1'b1, 512'hdcc948cfcd6f3cd3760d678a643ab0ff010000000095bdd5dd5c0b9579c7c6b0f3e921033117737e31acf8ab117b62ee54a25abdba306c71bb0c3d60097a332c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h047c4306f8d30e425ae70e0bee9e0b94faa4ef18a9c6d7f2c95de0fe6e2a3237, 256'h7a4d0d0a596bd9ea3fe9850e9c8c77322594344623c0b46ac2a8c95948aefd98},
  '{249, 1'b1, 512'hdfc50d9e551fd99c3ceeeadef83e2fab3f96000000003206a5e2b462805d83d6ef6280540f3bfbb229421d6f5f2794f117259f9dace4f82dd57889a74a0fcce9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h57d603a367e23af39c95dd418c0176da8b211d50b1be82bf5ef621a2640204f7, 256'h5dc3f285ad015c4d71157bd11e5b8df6a89e4b267393b08b5ad5013bdae544b1},
  '{250, 1'b1, 512'he4edde495afeff435a69e94a6493e4ec2c0b1b000000004c8e512f917698225b0189f732d3deb6d8c1c39b6b59e0701bd7f7605a521891358603454d151d8e7d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h11df6741021ec8cc567584aea16817c540859c4e5011551c00b097fcfc2337e5, 256'h668551919d43206ac0571fc5ad3ac0efb489bea599e7bf99fe4c7468d6c2c5e0},
  '{251, 1'b1, 512'hdf8f102f7c54ce2cb6ca609ce724818f7621cdc600000000c69bb15b7c33f6b27c75a153b581d47b99de18ccc8105fc3bb697f180112706c5ebfd6fc6c8a6322, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7451ffede471bd370406533436fc42a89daa0af4903d087cbc062fe7e54dbf70, 256'h590895398f22b48ce72cbf7c3d3ee1dd7fb0ee645edb0b1b1de35f370e5bf5ee},
  '{252, 1'b1, 512'h3e526c3c1f02aa2e007cecd9e02f7dc3d06f361a0c00000000f8e183a89a7218d8183a928d91c6bba47d950bf841396e5fedf9d87f66671deb8d2ebf63e39751, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hfc4c4d81da6f687a6426263193c1a680b67734a1b180647b8c76407cc4f0a9c6, 256'h56f775d372c9bee685374085be676c9cf31cf1f978a5e6ccb04e4a0761159cc7},
  '{253, 1'b1, 512'h7a750c1372a8d9b00991182aa031522b94a1a7f4509a00000000baafee68e65ef0a94f7983cfeb9241e0b7d8fd590a0d55b16041eaaabc38e982aaaaf6eb75e6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hfeb978ca33c46ffba47eb63bb40de7833e43d5654575b54de1fea3d1de3c8ad5, 256'h108078ba997bfa064521baf342c97b0c64bd25240c8fd0fd7533ae2d03081b70},
  '{254, 1'b1, 512'hb8df763eea0cf11e9945dc5667b0147cf8684d618abe1200000000917eeb543a4dddd7217ba71e998bb9c5fd62b57509b7cdb489bc3b64f66a70e4b5c12ffd2e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hcc61729698467ba53da199ff481fe7433f194fc96367907e8dc5e1d9f42b1e21, 256'h83dd9ef156e7c1f9c09b3bf86a4f1c88e5dd20cd74d997858e600797dbe74ad2},
  '{255, 1'b1, 512'h88670299bf6b255d331cd40c7154c438fab9fdd2b4319e440000000057a51b1cdea2812fd594a8cdd56b4f5cb069625524bd53a5f304653824d4afbf9bc58d02, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hd47f616303ff0eb813eac32e760ba30ad445e0af7dc57e70756104823f6a895f, 256'h047f2217b399c46a426b936a124980a6011f0896f51dbe07632828a72d7173f1},
  '{256, 1'b1, 512'h295422dc27dfac13c79d2028d3daed64c1dcaad525dbbf14a9000000003667b1baf41fd9137fa0bd8c3851590b206aefb6cde62fb4ecc23ae308e540e83a7f09, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hcff73dfa2bac67ce1340b25c885abb3e7979ef7f840f15d5f19e86640cdd40a3, 256'hc7d1210802796c4f251049ee08a2c29f5c71064033d17010c65bf2e94499381e},
  '{257, 1'b1, 512'h118422376e38638a08705cddcdd319e26fc8a2e6d4a4d1400fb70000000005687b339ec07f51592f6e254c9b7291fa2d0302df9fb2702857e3f69bd4fba01654, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h10acaf9c485ab1220355b95be269f124e12eb252f2224b0fc50785eb2ee3df45, 256'h32443b557efc6896347fa778e1fcf33cbb769c9a7da896b20d93fea7c2791ea4},
  '{258, 1'b1, 512'h5a4801a1f7ef2afbf8e0e76cbd6e07212568cb47638e22e55f8e6c000000003a2aff81ce04258211030942fca855cbc0ef482027b17a7ee523b15483afd91355, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hf919da0651abc2bff994a879d2778fa5195d57400e003e8dd6adb3fc7a0cc4cc, 256'h9b945d06bd119665b278a59bd24fdd2350817d0be87997bee57b70c479d64a2d},
  '{259, 1'b1, 512'h057d7524efbce651b92e0a70e4454156e7cd4b696c197c6a064032c100000000768565d4af2019fe3247dba91948292af777f107fdc9c3b47659eaeab26ead77, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hcc38e7a018f6d70b2d9b49120cc9b4a169f2f72238821a86b81f553b6225d24e, 256'h276efd8bf06ccce07c7aae35eaac3bd1c374dcf0cf0588d5e0e4171936688636},
  '{260, 1'b1, 512'h31ccd924b687a2a6b70f4888ea911ea38a686e56e5540ea692ca3174bb00000000246ac69c46506bd8fe924eec33b33ebc9f508d4251c459fdcee3b4c84d4ea3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hff85ad66621991c318b85cef73c576cb2a8d43c568c1aafc85b40ef2a9a6b41c, 256'h732a79e6837ebf8434fea6e7fefa948f506ae455c1a3eb36a030185a23037d96},
  '{261, 1'b1, 512'hc7b70cc4a55d55342487a4469ad2243ef6d6b69f11604b8c12baa03dd3e10000000014df0db29a9d4d54b26f4047f3e0c739f7a260768b20589254e1235fc590, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h33f016e51eef9b1136380cb8b84c6b38b107e24c6731bd07cb1c7f4a29f33a83, 256'h36b177bb8be94c8be67ff3a41fcc4d22b5c9eb377da713eb014ae01c64ca6dd7},
  '{262, 1'b1, 512'h1634df8a3271a99f360e3bbdcf789d24bf4bb03e3114ee9f0fa930541f1ae0000000008d976fb74f27eb316ce3a24d92a53833e600c353300f5c4fec6b28c581, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h929413ee91f27454d74e91370a10a86fc98ac7305c8ab4ca59752bda3a7bfc37, 256'h483b47a26a0d7d2e6bd37d351d9ee37c5ec2a4686d884d78b6beb7f6b08c50f9},
  '{263, 1'b1, 512'h8f90b6a8ecbb870dc24832b1f4719aae2d8eedd7faf97848b08d2b528abf5f44000000008877a6157344e6a9dc43b90c8e2dd7ab9bdc5237c912e094660d0878, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h578202c7d0abac93ca43dde3cb44414e5601c1eb557604cb9adb4bde0a12633b, 256'hfb9a7412e307aee95ef4b53540571a21559414e5306794ab5182cfb229dab3e9},
  '{264, 1'b1, 512'hc0891fc626ef4b106fc00f5c067253f26a2868d09aa2ce029466f353ba525e757100000000a3cee37421995445fae741697659a406394c870d8bdda130080d15, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h46d45ad0bb75b8639d0e91d8450fc31887c211328a5784fc83b4cb7f5b962c1b, 256'hd6751d13ede2079b7aa1d822bdb32d7f3cf00273a1ff03df90c0ec7c62a47568},
  '{265, 1'b1, 512'h76527097fb3945436a30cca60392c170abb7ddf6ddae93e3ff7651d468eb3e14865700000000bd314c31706f8e4d1d853b151f5afe680e13cf2f255b2bb697bb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'habe84c941783d5ced284fea56341ecc68d6bdd3196d318fbd074641f8c885bd5, 256'hbdea3c44d48e01aa40935c1c9723ff733199563440f26b4ecf0b444b0418d9f5},
  '{266, 1'b1, 512'h41d43cb27d4db522756dd682826eee8d0f60163c7f3ce67a39d89d7d89e24818c354ef00000000cab56830cd18f7bb9a7d1b2440fde06ce647518fada2dc988a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h05277cdbf491e336fe81be24e393a161a4fb89112c9ffed1ee6649c406713408, 256'hab6934332e68e108bb0484d21c457dcf381a620c3a4712fdbfeb658a3fafd60c},
  '{267, 1'b1, 512'hd34ac40ed5ab79a4e5ac1e4081e0e47e4fdedac1555b01ab62a13ac0ae9dbc3c23f799510000000010116f328ad1db0cd68cd1db9e1b34b5a52ebe9b8e372b78, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h293825737c8c14430ed10dbadd7da337275f9b61d1d26377f778ffaa00c139de, 256'hcdddec267a8678c96829bf6c1d6f38322e119937cfd2fee01e9dc9525f43ed6b},
  '{268, 1'b1, 512'h8b5db6db13b1f5e609965dc38215d14ccddf66a9d86505a67cca37f13cc420803c1df80f4700000000b044bda09a83e4331aaff90c4faceea315e467f5fd91d4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2041fdd6111c45dfd29e750e082dcdadc9a584a8a2be46580fb0ba3b3dc65862, 256'h421824fe987e4172a0f8bbcb7bcd9e1b073b7742ed9f9df98f2a1a37cd374ce3},
  '{269, 1'b1, 512'hc771e022bc376ffbe1f513bcff11884e790e53878c197014931f6360c517ce8de1c059d091cf000000003c560cc443a6f005ea58917a52ca9bf60163afb16ce8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h267941db660e046ab14e795669e002b852f7788447c53ebef46a2056978b5574, 256'hd00183bcaf75bc11e37653f952f6a6537151c3aa0a1b9e4e41b004a29185395b},
  '{270, 1'b1, 512'hd9cb55a3f1ec161bf6caf0452bd6d6c876b35dd1000eefe18378afaef6280348fd799e624e573a00000000085b3b24635f5c10770090ea935f198728655e236d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5dcd7f6814739d47f80a363b9414e6cbfb5f0846223888510abd5b3903d7ae09, 256'h43418f138bb3c857c0ad750ca8389ebcf3719cb389634ac54a91de9f18fd7238},
  '{271, 1'b1, 512'h0caacc1f43ee27ec7ad5269155a66172ac310d4e202a9b7d3defcfb07ea8da85415ac2b116e665830000000009887d6c7da6cda824528345e14a6675de23988a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5e0e8cc0280409a0ce252da02b2424d2de3a52b406c3778932dbc60cb86c3567, 256'h93d25e929c5b00e950d89585ec6c01b6589ae0ec0af8a79c04df9e5b27b58bc5},
  '{272, 1'b1, 512'h5d761de2a231df86c0fdd90da20e5811f7bd9bebb3f1966359b8fdf554f79f0bdd32ca06410e70e61100000000ed3d4140a60908e85f7fcbd26dc792bedacbfa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4fcf9c9d9ffbf4e0b98268c087071bffe0673bb8dcb32aa667f8a639c364ea47, 256'h820db0730bee8227fc831643fcb8e2ef9c0f7059ce42da45cf74828effa8d772},
  '{273, 1'b1, 512'h78adfad2734b7baf32f4e0201bd6c3e9f6c1763cbe35858a0f56466db34dd98a0fbf5b2a71afbcdeebd400000000d3da1a5035406b39aa13c126a3946b6c6a5e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hc60cd2e08248d58d1639b123633643c63f89aff611f998937ccb08c9113bcdca, 256'hac4bb470ce0164616dada7a173364ed3f9d16fd32c686136f904c99266fda17e},
  '{274, 1'b1, 512'hf1d6ef224f72b83a109944afbfb34ae1f70d6e50eee54a91faf8ba0fc062563113d988f2b826c055ecc61e00000000554878a7e761e75fdf1ed2ad2d138b2974, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7cfdaf6f22c1c7668d7b6f56f8a7be3fdeeb17a7863539555bbfa899dd70c5f1, 256'hcee151adc71e68483b95a7857a862ae0c5a6eee478d93d40ccc7d40a31dcbd90},
  '{275, 1'b1, 512'hb33f308c5b107050cb2e513fabf8b896e52c85852fbe32308bee8b8661121bdac78f52f924cf3d5690ac92d5000000004f0f619e72ec1464166078ba3f508a66, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2270be7ee033a706b59746eab34816be7e15c8784061d5281060707a0abe0a7d, 256'h56a163341ee95e7e3c04294a57f5f7d24bf3c3c6f13ef2f161077c47bd27665d},
  '{276, 1'b1, 512'h0392f8c2dc961605c5693d9452731b6a8292ff57d6995aeca0dad3117459668ec7809dc09cf154170fcd624be50000000026e3d92dfdf1a2abd09392468117c9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h16b5d2bfcaba21167a69f7433d0c476b21ded37d84dc74ca401a3ecddb2752a8, 256'h62852cf97d89adfb0ebbe6f398ee641bfea8a2271580aac8a3d8326d8c6e0ef9},
  '{277, 1'b1, 512'h9dda0539bfe47c75bc00b014dc6046c9db5d7a5723acddaccaf2aac7a9250b732a80cd948409f132d1dd65cfe91600000000d53c76be9f75fc6927f818acdaf7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hd907eefa664115848b90c3d5baa0236f08eafaf81c0d52bb9d0f8acb57490847, 256'hfd91bc45a76e31cdc58c4bfb3df27f6470d20b19f0fba6a77b6c8846650ed8a6},
  '{278, 1'b1, 512'h572e1d736d78c42eed5ffabdfb25b5c7908aa60728ddb3d36a24c285db9ab996433827aca9e23716c3baabbbb4527600000000b9c1a728fdb6f65c10935e9514, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h048337b34f427e8774b3bf7c8ff4b1ae65d132ac8af94829bb2d32944579bb31, 256'hbd6f8eab82213ccf80764644204bb6bf16c668729cdd31dd8596286c15686e8e},
  '{279, 1'b1, 512'h81b675425e8c528a0a51b23413c8b796411a01b207e0bafc5bd2a46b05237be84abdae1ebd492fca053bf7e3133392720000000086ce63108f1dc5a3b34c575d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hb2bc46b7c44293557ab7ebeb0264924277193f87a25d94c924df1518ba7c7260, 256'habf1f6238ff696aaafaf4f0cbbe152c3d771c5bfc43f36d7e5f5235819d02c1a},
  '{280, 1'b1, 512'h11c203ef3c8978266a73147233f7c9c9d16108a07847ff587f1e865f28519e7a161664edb56d9e791fba0717124717b3c90000000013c59e26ab63c4a99b871c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h40d4b38a61232e654ffd08b91e18609851f4189f7bf8a425ad59d9cbb1b54c99, 256'h9e775a7bd0d934c3ed886037f5d3b356f60eda41191690566e99677d7aaf64f3},
  '{281, 1'b1, 512'h5de83c97136ff31a90ea5053ff256d522819626ae3734c460ea7681fbd0a94538ed840f3bfbf8055756e761d8149786b8cb000000000f37f36e4d32d46cb9bd1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hac8f64d7df8d9fea005744e3ac4af70aa3a38e5a0f3d069d85806a4f29710339, 256'hc014e96decfef3857cc174f2c46ad0882bef0c4c8a17ce09441961e4ae8d2df3},
  '{282, 1'b1, 512'h4a5e1e8c073ecb2832fe0d0df42a72ce225ea97ce093ed320aaba00cab25ec3e90a6aefaae72ad40273d7309e40582f40a37c1000000000b1e8576da0eda555b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h41b3766f41a673a01e2c0cab5ceedbcec8d82530a393f884d72aa4e6685dea0a, 256'h073a55dca2da577cafb40e12dd20bf8529a13a6acdf9a1c7d4b2048d60876cb3},
  '{283, 1'b1, 512'h9f920bb92b4527d54ff6877b80c81585dc4d3d1e96fce780b030f9f371f8a1b68e2e7a86536acc3ce96737bd5fba0ff669f6b1600000000000b5868a36cfe6c5, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1942755aa8128382cd8e35a4350c22cc45ba5704d99e8a240970df11956ad866, 256'hf64cf1e0816cf7ac5044f73ba938e142ef3305cb09becb80a0a5b9ad7ba3eb07},
  '{284, 1'b1, 512'h99f941e73ab790b224ce0a799133f6b04eb9bcfb2fd0ec84b8e7d5dca6ca50d2b1ae4d31c57e2e54f97f59b6a10d0758cfb3e46500000000909d4fabd9d1962a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h51aba4ff1c7ddf17e0632ab71684d8de6dc700219ef346cb28ce9dafc3565b3b, 256'hb6aaebe1af0ad01f07a68bf1cf57f9d6040b43c14b7eb8238542760e32ce3b0c},
  '{285, 1'b1, 512'h202e258cee0bca789ccd4c29f3835362b6f1f53faded0f1d58f4ff768f6202a6de3ee3b922546127fecfdf1c0446605751df9b7fbb000000001a8a11a3e383f3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h91efbfcc731650e9f004c38b71db146c17bf871c82c4e87716f7ff2f7f9e51d0, 256'h089ea631a7c5f05311c521d21ba798b5174881f0fd8095fb3a77515913efb6e0},
  '{286, 1'b1, 512'h8c4a184638926ecd8f6ae279181f9171181295757e3eae5b5a0de2fc0281358973a355e4820da4ce0c69db549c72ea007f80ae990565000000009e51983c039c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4a7e47bd281ea09b9e3a32934c7a969e1f788f978b41585989f4689e804663fb, 256'he65f6bd702403cbbed7f8ad0045f331d4a96fbf8c43f71f11615b7d1b9153b7f},
  '{287, 1'b1, 512'h92eabef5ab4296dba863345a2f11c2bc8d32bc02731323a19a88897aa1421f384448516975b6397a8e627fd3cb5a5dd6ee3c50226b18860000000077b18d5c83, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hc795f5da86e10a604d4f94bf7cac381c73edad1461d66929e53aa57ca294e89f, 256'hbae784ab6c7b58332ee05e7d54169edf55ce45f030e71ae8df63969fb327a10c},
  '{288, 1'b1, 512'h4cb05f07197bd719557dcfbe1edff395550b275100cb073ecb4a0987621f83a5f041996f63fececb77a30cccc5f8067e36f650f7defb611b000000006a949e2d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hea68b24843b225f505e01c0e608b20b4d93e8faf6b9cf70cf8f9134a80e7b668, 256'ha3abc044b4728f80fe414bdc66f032b262356720547bec7729fad94151c6adc7},
  '{289, 1'b1, 512'he744eaf4e9c4c17549ca3907721df98de95b69d07d56eef509d4740a3cb142bc61b6c4d108676526d5a77188977d924dc9a8adf6c01adc35d6000000007f3077, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hbfe7502140c57a24a77edc3d9b3c4bc11d21bdb0b196977b7f2b13ac973ad697, 256'h947a01da9731849d72b67ef7bc40b012480fd389895aad1f6b1cdbeab3b93b8d},
  '{290, 1'b1, 512'h4fbf285c9be6083627ef151df0d2c5fb00b6edcfc44216a30467a4fe268214ab66dd9be898bea57b48f6499d09d4beddb7c9e8bd813fe7c1cacb0000000054f2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3434ee1142740a0ab8623b97fc8dc2567eda45dadf6039b45c448819e840cf30, 256'h3c0fac0487841997202c29f3bf2df540b115b29dc619160d52203d4a1fd4b9f7},
  '{291, 1'b1, 512'he698cebca57a541614e179f28ba51cf82fa0fb4300f81df5fe22b635eb4441b496a36ad280999f503edded3ae1cab1700758b5ae80ce33dbf25c7300000000e9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5338500e23ba96a0adc6ef84932e25fbad7435d9f70eb7f476c6912de12e33c8, 256'ha002f5583ea8c0d7fb17136d0ee0415acf629879ce6b01ac52e3ecd7772a3704},
  '{292, 1'b1, 512'h43f5ecee4c9b5bcf2497d9753beb1eca8a01c143f8b50518e83bc7f3f62d049b03430a6dbc9236d54b7ef5475a232e3de9160e9649e3c8f46d2f1f7900000000, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4ff2d4e31f4180de6901d2d20341d12387c9c55f4cf003a742f049b84af6fe05, 256'h0312f38771414555fa5ed2817dcc629a8c7cf69d306300e87bc167278ec3ef37},
  '{293, 1'b1, 512'hffffffff4fbe152fff953f198736b155220dfe633b6fc7aa5bb392cb96cde9fc658b17828d0d04ece0f6e35ed6bbf357b86665cac7735a3b9c85c038d4a85019, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h51d665bad5f2d6306c6bbfe1f27555887670061d4df36ec9f4ce6cdfaf9ea7ac, 256'h2905e43f6207ee93df35a2e9fb9bc8098c448ae98a14e4ad1ebaea5d56b6e493},
  '{294, 1'b1, 512'h47ffffffffa19c2322e79638701c393ec0df74b5d27fb9ea7cc3e3dc8badffcac83dd8c409a22c2d7a64b5693f153f60264487aabe5df546115cf2eaae415ac0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hb804e0235f135aba7b7531b6831f26cc9fb77d3f83854957431be20706b81369, 256'h9d317fd08e4e0467617db819cde1d7d4d74da489b2bce4db055ea01eccfafcf2},
  '{295, 1'b1, 512'h391dffffffff5a981c0576acae266e7b35ecdfeddfeb6db903e9f4eab200dba039b146517f0c5b418d096addeab6d0962a6f77c2a2a552748b788c07796553e5, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h8ab50ef3660ccb6af34c78e795ded6b256ffca5c94f249f3d907fb65235ef680, 256'h49d5aaeae5a6d0c15b286e428b5e720cf37a822ede445baa143ffae69aba91b8},
  '{296, 1'b1, 512'h8c8ed3ffffffffd5bc0cf4859c831b89860c28ba17ff5a259b6982325be66498c4ac3119da331db0976678878c73473aec528a7107d0d9b1a17dacb9a9237b1f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h571b9c46a47c5cc53a574c196c3fb07f3510c0f4443b9f2fe781252c24d343de, 256'h68a9aebd50ff165c89b5b9cb6c1754191958f360b4d2851a481a3e1106ee7809},
  '{297, 1'b1, 512'h531341a3ffffffff263c81971e877fd7cd8308b0d536d7fa3c88e3beaad332ef664f76387e4c43dee6c0a06423b18d1b1772f65acb4f9b672b97a648cdd25929, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4cb7817b04dc73be60d3711803bc10687a6e3f4ab79c4c1a4e9d63a73174d4eb, 256'hce398d2d6602d2af58a64042f830bf774aee18209d6fb5c743b6a6e437826b98},
  '{298, 1'b1, 512'h2639a8ec01ffffffffb54d98af88ba2ae383d69bee2f5fadda599d58796fc766130e3fb8f4ec1afceb8a1c1faa3ad305a0fdd65796adf8ac579c1306d5f0195d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h684399c6cd6ebb1c5d5efb0d78dce40ebd48d9d944eb6548c9ce68d7fdc82229, 256'hcf25c8e427fae359bfe60fa02964f4c9b8d6db54612e05c78c341f0a8c52d0b5},
  '{299, 1'b1, 512'hd9753a5a8b1dffffffffcac9aa24c9d687a2088ed837789e72d457d0bc67f54860087c3f0509744e0b461f88893e2de6c757705670006c9e9e8c4c3757fcb160, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h20b7b36d5bc76fa182ca27152a99a956e6a0880000694296e31af98a7312d04b, 256'heeeabc5521f9856e920eb7d29ed7e4042f178ff706dff8eeb24b429e3b63402a},
  '{300, 1'b1, 512'h9a6bf9edc61a22ffffffff703f4706318ef947658ec44c90cc1630c916924f1635efd88bcb900db41dad160ea33f8176397bb8593e19199207ca7d57bbd28305, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6b65c95e8e121d2e6ee506cfd62cb88e0bfb3589da40876898ef66c43982aca9, 256'h09642c05ad619b4402fd297eb57e29cca5c2eb6823931ba82de32d7c652ba73e},
  '{301, 1'b1, 512'h4c18a4947b15af08ffffffffb9de1de3873b4c26280b1286a51715dcfd1242208ad49b2aad0864d5a4529e4a653d7a6355b7c1747fa9d876159d43806661395e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h67c74cbf5ea4b777bf521ace099f4f094d8f58900e15e67e1b4bd399056629ed, 256'h3d2884655c49b8b5f64e802a054e7bf09b0fc80ca18ebf927b82e58bb4a00400},
  '{302, 1'b1, 512'h6e50953fea8dfead2fffffffff824e02147d010595358c98ec376055cb9ddc1dfe6d3874cf38e8a98ef0664fd3b10605bc14506eb7e46460c9db81b10e2f6730, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h79a5e40da5cf34c4c39adf7dfc5d454995a250314ebd212b5c8e3f4e6f875feb, 256'hb268920e403ba17828ff271938a6558a5b2dd000229f8edb4a9d9f9b6ac1b472},
  '{303, 1'b1, 512'h1539fd34220ed16ae0b8ffffffff88a04bebde47a3a94f1b86bc687c2ce7648caa7d42ac8693b5704e401b7c9f4864bbafe3bcf761d862739eaee02516a0d707, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hc8b13006c3a51a322fff9321761b01de134f526be582b22e19693c443fc9fe46, 256'h34e7f60179c6162ab980fcd58f173b0e6c30b524d35c67921677522dcef843a1},
  '{304, 1'b1, 512'h69e3c78c7125bdee7184d6ffffffff274929ae7dcfc4692b84880a518de1790a758005ef7d4e29377cd891eb08e9fda55ac99a11b4dc9a15ceaf8887ae941fd7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3513db745489a487c88a6cedf8795b640f8f71578397bdabd6cc586c25bd66ad, 256'h99a72cd3f0ca6c799149283ca0af37f86b88200d0c905bd3c9f1b859e55b1659},
  '{305, 1'b1, 512'hc3b630a45b21b937bf78ef4affffffffad33da42317364a1090ed4446da7738caefc807ed99c92f85a6f6ba946f99284d4b9793896bc5e0b6f93cf1b09b35a6d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3a6386afb08f7ff8140b5a270f764e8706ef2830fb177446f7b4eeb8a25aac64, 256'h4b70854b38c29245b2b980eba10ea936c68a38c1da5255ce2386db23afc7c06a},
  '{306, 1'b1, 512'h14f3b0fc1795c9d400d904ea0affffffffeabaaa40c2f532e33f6c61620d23188712a838f9bd1502b2a5c321117ed6007ccb48b375c581fadf340b0d7edcac93, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hb8fc54a8a6be3c55e99c06f99ccdcce7af5c18a3c5829726a870cc1068458f64, 256'hcc7237c39c8e6a4a1c8c62f5f88636549c7410798b89684c502c3adfe5fb7ad2},
  '{307, 1'b1, 512'h386b3f08bc91c7e18354f3d46de4ffffffffbf492f2bf174abad52337a99f29dda6891d96f85efb667480bcad7d2482ef7f32a314b4dd39576ef560bf01fefa0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h47b460851e5607f2021626635c565a63f78f558795e1b330d09115970dbbb8ab, 256'ha6a9f4f213e08d3c736d3e1c44a35140cb107619f265a5b13608ed729fd6d894},
  '{308, 1'b1, 512'hcd86d593a60faa34608d5bcdb2e878fffffffff06003c116f812eecd35fc6f3cccc1dee24c5cb89cfe9d41b0defa4e5d16b1d9aa4897e6efc838a8a6dd5f22aa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h8cfda4f7a65864ebbea3144863da9b075c07b5b42cb4569643ddfd70dd753b19, 256'h595784b1ab217874b82b9585521f8090b9f6322884ab7a620464f51cf846c5b7},
  '{309, 1'b1, 512'h7939a3e06bee091634b535adc98afd56ffffffffeb0206c5b2cf892d2c8fbb5a2e105567cdc4447b476525488611a085b870e498a13b891cfb9a66ad725273af, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4cd6a45bd7c8bf0edbdf073dbf1f746234cbbca31ec20b526b077c9f480096e7, 256'h7cf97ae0d33f50b73a5d7adf8aa4eeeb6ff10f89a8794efe1d874e23299c1b3d},
  '{310, 1'b1, 512'h180c134c29d50916f2c3b32bf43382eeb0ffffffff6178b5edf0856813b75ccbb537c57758d3e55c190bd8e648a79c5bc6a62e45f2f037aeace1733bb7260707, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2e233f4df8ffebeaec64842b23cce161c80d303b016eca562429b227ae2b58ec, 256'h46b6b56adec82f82b54daa6a5fca286740a1704828052072a5f0bc8c7b884242},
  '{311, 1'b1, 512'hf2694ba9c9a0d83faff7ff2f06f0495682e8ffffffff1d5cf19e626efbbb1425dd286e93044edf262236a46a82638145b4d15c18aa6e1edc919e22bff3a9c5aa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h549f658d4a3f98233a2c93bd5b1a52d64af10815ae60becb4139cac822b579c3, 256'h27bdddf0dbcf374a2aec8accc47a8ac897f8d1823dda8eb2052590970b39ce2a},
  '{312, 1'b1, 512'haa2db4394e6e52a9f0485ea08186ed648a109affffffff19fae34ae6524a6abf956c07617b15896bd3dff11cdaed4f9a2769cb4dad0b0e007b66c06fda3f256b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h9fabcc1e5fd965226902f594559e231369e584453974e74f49d7d762e134fb9d, 256'h293cccc510793bac45ce5da2bb6c9e906437f59435ca206655f74b625df07c7c},
  '{313, 1'b1, 512'h59ce78a87d80e90e1e6b70def3179e12e78cd5f0ffffffff11eee1f43a7030f096c301beb60d1fc2be04d27aaec7c385fb9aadcd6fa37cbea40783569080dffd, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2e5c140fd6f5f823addc8088ffaae967e7f4897274316769561dfb31435825d9, 256'heda47327d7cfae1daa344ff5582a467bd18eb9f01caeab9c6da3c0cc89df6713},
  '{314, 1'b1, 512'h5d07345f237708f45b49a7286977f331a27c8cc58bffffffff492a29a714f16596215046376e8d35cebaaa06b73f14ec0731a0607ab89c4edee5ad7f575c93af, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4c11e3b7efbe3908ad2118e54d7d34d6c6eb4570bf7fdb11a7679fe93afa254c, 256'h712e90f421836e542dac49d10bb39db4a98b2735b6336d8a3c392f3b90e60bbe},
  '{315, 1'b1, 512'ha6d55690f7fe8dc6a67ac00e5f136dab1f6855b53643ffffffff2585eedbf8e7c3db326f7fed8c48851376d7b1a34dfd79aa6837d19b05becbe8b8d122d1baf7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdfb4619303f4ff689563d2275069fac44d63ea3c3b18f4fb1ac805d7df3d12ec, 256'h68e37b846583901db256329f9cf64f40c416fba50dcb9be333a3e29c76ae32db},
  '{316, 1'b1, 512'hd42f5eb7f42a9dd25a5d9513de8b6ccd5bbbd029263799ffffffff3baff5bcc111d8fb4f14fc4aac37a1dc5633df840644aeb69aa87f390c090e6730bade402c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'he70e8e17bd758ff0c48f91cb2c53d293f0f5ae82eb9dfe76ab98f9b064278635, 256'h21dde32cb0389cad7bdf676d9b9b7d25bb034ad25a55ea71ee7ee26a18359dd2},
  '{317, 1'b1, 512'hbf0fafaf135ee4e03b991ef87e6e9377150ae255e043de57ffffffff10002deb92f4bf4c1770933d3137b0165ebcf81c8c3387c21457e0fe0c39c7c7947837b9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h421397ecae30617a5a6081ad1badf6ce9d9d4cb2afdabf1f900e7fdb7fb0af5a, 256'h57ca89dc22801c75fdbefdaeca65c675625f94de7d635062b08ed308df5762cc},
  '{318, 1'b1, 512'he0dff3b5ebca4c971f1da5a6726d24519e4ca71f45a548d85fffffffff415d9ea4bcfbe4749c275d6594e8ca8b76166fc90eaf2d9f466b0f0a5ed8c14eef030b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0610c08076909bb722fba105c23eac8f66b4db1d58f66a882fc90d59acdec8e0, 256'haf59e8d570761cac589d49f11c884007f7ac1eea1a44c6f3fdad1d542187d25e},
  '{319, 1'b1, 512'hd9a9dae1785ef8a49d7c81b0637471693412a29484ea1cc780d5ffffffffb70ab50279ba56f6576dd87ea0cc08ed51afd395238936b4aef7284700c8d5aa9f05, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h59a1181cab0ee8ce94ab2b5ab4f4b13a422e38efe69f634bf947485a5b9ea49c, 256'h9b3c913d98a4ab15f6a39f1802b8f2d28559aa1f8d03a3a88df00c89dc293a97},
  '{320, 1'b1, 512'h75c7b98cfddf04426dda027ad897cd5ba9d5318c27288ec0f6fb67ffffffffb744ccbcda470681f3689c70425ce514d035e05dd133da5c2a104980f4ffb91014, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h8cae6c4dfbf901bd66ab82541011fa15c8e90e2c18c01bd881acaa2b63cb587b, 256'ha86acf943f29cef91d1b66a7de5547df6cdfc45dd7bef816dcb8de9f5a425d2d},
  '{321, 1'b1, 512'hccfcfe85e6d12e377ff1bec515ce149719d86cf3591b3dd8d4344022ffffffff60380790c2be6a944f31e63ee7b421a42ec5ab43f84f05aadc5ae5c42a6455b9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h8b00c74b86474d782eac9974aea606d8f7ee78c79597e15687021f5991e86acd, 256'h309dfe3686648eae104e87b3e9b5616a3ad479ca4f0b558ae4f1e5ab3115346a},
  '{322, 1'b1, 512'hc445da85686a33c8af5997da14f197df87bc3ff9f277b46831c87f8147ffffffff0970446a79a2c801e1a6f9c03509ae9b782a31b3b15dec03f5789a8345e14a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h433a915504c977809634a36fcf4480e4c8069fc127d201d30dfdb1f423c95fd4, 256'hbcb1b89aafd50a1766b09741fc6a9a96e744ae9826d839bf85ffb50a91981773},
  '{323, 1'b1, 512'h6a94c0cd0809f1ee1c23039f735f24a0a006a0504c295289507a9dc93e34ffffffffd7127f6a21cd1ec975e05b1a8d78144da6293f4440723e7d6062dae06a1b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4b69abd2b39840a545cdd4a72d384234580e2fd938b7091d0ecdb562780857db, 256'hfdab9957119e0a4092af82f6cc29f3c8a692671ec86efb0a03c1112a0a1e0467},
  '{324, 1'b1, 512'h31599cefc10a3c6d549bab5b19bb49d01fad30283d27c8a4905d18cf61e045fffffffff3efa7e2362af0fc827c4bf245dcd58374b350097d26ac996598012290, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdab9d3686c28363ad017b4a2b36d35bf2eb80633613d44deb9501d42a3efbd38, 256'h1392a562d79f9ab19014e4f7e2f2668259f3720a76c120d4a3c3964e880f7679},
  '{325, 1'b1, 512'hefe7f8f35a94b65eb3a9299658db8b8256f29f2df969035fe5769c11e85c9b7bffffffff61e57fc3e05c9a1eaf760ce1b13dc6ddc5516048677e1fcd420a6427, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h23f94e47b440ce379b74c9311232b19a64e3e7c9b90da34b0c1c3f3d7af28105, 256'he1425903b1479c2ce18b108a6d1ec8b7a4f0f657dedb00de3a3ceea7fdeee9be},
  '{326, 1'b1, 512'hc5c3daa9bce3e7422af1de2fdc992b34f5c8ef3fd448b45f2426e1677feaa86aa3ffffffff6e9d87ba471035c9beb5d2c94f3bb0dfb4c48298a8615840c621a6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h9d706a8fa85d15bd0c3492c6672dfe529f4073b217b3947b5b2cfd61f87ccb71, 256'h6aaaaf369f82a0e542f72ded7d7eb90c8314ffa613a0ea81da1c8393dbae2bac},
  '{327, 1'b1, 512'he36dcaffe4916e59e41b560c2961fba82290150d1b262323c674311ef6c87564c8aaffffffff573ce47a2b2f25bd4f6468ef2788ede75cd3b7293ad2bdb46617, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hac77918c4085c8a7ce5020b00c315629aee053a445cb4661eb50f6b62a47da29, 256'hdf2aea2b9c11a6ce39d3cd9e1faf4a53057e0b1b2e48a324be9e773203fe9fbb},
  '{328, 1'b1, 512'h3f4f00f697d80c258cbcaaeea0f4fa499e0675441a078d32627378ae08c27dc9e8b60bffffffff59976ce86a303743b716e53422d7a17166a185fac1b7722d2f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h9db2dbd2935f147fae7f6a95c8e2307bd8537c3d96eb732ad6d5ebdd89bc754e, 256'h93a9ab99d2de9d08fe0a61e26c8fe1ebbf88726e4b69d551b57d15f0ae16df5a},
  '{329, 1'b1, 512'h21b10973b98ea1dfd2b0d7bfe4adf9d4e8616759177daeef38d7aef0d95d226ec8e1da39ffffffff43f8e40342757a93e72541afd7a58ea2205891c13c72a8e4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h769f70093939afbd1fa15873decfa803ca523ace8040280ba78cf833497722bc, 256'h369875aba5e1ced5a4ca8444ec9399a38038b00e153a0ae34d9b3c9781447eea},
  '{330, 1'b1, 512'h3be3c1c0f8b8f6b9c476455ceee9edbf99283f1eab4a28ace9494eae8da166e4aa1d5def8affffffff3d69a06db8c19c0984bdd10df6ede19e4214183d3b0762, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h26e5182b9822550ad52f46ad80781d6bef3d110a204db5e58a0746f796982200, 256'ha9418e76029ced0cf78a571a9e59ad04086e91f70e6813981bb33c1dee891165},
  '{331, 1'b1, 512'h14a2049293367e5ace79214bfae58e1007b4977ba9dbd787dd703160651e580fc6de8759ef1affffffff483224ed924c7a2906cccf6b3b39e1af044f2a7047fa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'he7bd6aefcf7b27e1f3fadbe713f9adb3d23398e88200cd2e94989c9d12e92177, 256'h9583e0de3b76f8d4b1e634a81cbc34af54e2f8599f3684ce48d372760c8204c4},
  '{332, 1'b1, 512'h745beae01e0b877f882a42a6339b12080d956dfd5fa03fc87f6c99096ae69833fab59c416b092afffffffff5deea8d387d1ecabbcedd6c2334cf7eaa7aa55d84, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h8638ed7eaa83609a01a6af9c52ec9bfddda90442b1e6031d61cfa22e48b2e1e2, 256'h20c284d596f71c6c8df732f5a5a2006302301e1a792e2b39663d93a9760762d2},
  '{333, 1'b1, 512'hc09dc1025bb9bfa3ef093eb420b7712374f3164db871d4cb44b8ebbeec2d5b415a73427419c5e399ffffffffb45643293f60ae63fb9ff87c56cb45252c8c7c29, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h61d924307a96180b06383608ba91674e15c3ea06ff2534412b93a587dde649c1, 256'h59b84aa2115b2547edac88088ca6313e9fbe1ca6a361c7e57938f9dde3f4349c},
  '{334, 1'b1, 512'h5f9b29b201a8f63acd7387dd71844b5ee67ca50c5a76a2b273a80d167abbdb6727992779f49b848976fffffffff2d0eab3e1c8f8be0d76338c7e8c92174b32c9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h424fcfc3fd63d128c2eb125e88c7fe5d283b63470a786b82783edbb8a0b7a6d7, 256'hb11548c2cd7fce9d44e795ca51af0b2f6a5180e9c9be0314007ed9e7f4bbe5e9},
  '{335, 1'b1, 512'ha76f6918ab70eb9171fdaecc8add5917f130dafbb7077543007be1aa2cd3e446114f1fed5989c6275e0fffffffffd7f5a47bd23e9cd47f4572a1d1146b38972f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'ha5f747ae6290fa9582c6ce8d5608621d495f061551bc4531bacba586a563b184, 256'h62faf8f92291e12812835b3f1d43c967bceb885b110bd06e5a68e2d74781ae2b},
  '{336, 1'b1, 512'h1694c34168745c74ab9fe8224e6058e045c73458f7e43e3884e3ed466f716a7406be99e0ef57710a1cac21ffffffffd497d0337e572f1afbc8b6b4f41a873e22, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hb731dc0d92c2cc7a605d78233f7814699bdf1cab2df297b6844eec4015af8ea0, 256'h39b1a0cc88eb85bcdc356b3620c51f1298c60aec5306b107e900ffdba049dd6f},
  '{337, 1'b1, 512'h3c28cf3e9527af87b483e6261fe32cee8e67cbc04b983566b27f8419a932186bce21c021eb58c8ecb0b707d9ffffffff035e36909fbfd832447041be74d2ab4d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hef73c4fa322da39fb6503bab6b66b64d241056afbcd6908f84b61ccbbe890433, 256'hf1ef85413e5764aa58a3128ccfcf388324fe5340e5edf8d0135ae76786ce415b},
  '{338, 1'b1, 512'hea6682cf1dadc5f218d6530a15452aaee8857a4318ef3da3cab58358a2e5d0f8fde22dc704453fb8056d224426ffffffff4335e1ab7e6e6c5f3b0a789528694e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h694cd30e2ad0182579331474b271ee2d48723bc8415dc6513873586ce705b76b, 256'hc5ac0c0ed5a4017d110cb45d63aa955dc7dc5ce23e7965c5397c3ff46a884636},
  '{339, 1'b1, 512'h0477828c9cc5710ded82ab21dfa5887f29edfb47548a5a99ff8315da76be5f67922c0a5de1cb7448a3a79b214889ffffffff7dc823ffb5d2fbcda33e63489df0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hf38b2236be3024e10b894ffb1cc68d0bb8d4cf0fcd2cfc1779f8883765d3cd96, 256'hda69cd0b74c25566d60a486edd559fc39d569fb2751445a4798df8a36891802c},
  '{340, 1'b1, 512'h17dfd1c9bfab4afc7d5ac126157041f4c4ca4a04aaf17c45e47857c384fb415e4362041ec3e91609325b7e4c9fb1a3ffffffff9d3efaa9406e392a0dea1ea309, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'ha881732c205a0b4b95669c00756fd91973450109a46f17d5a9d971b5e92b9aa4, 256'h8acefdca4e06c16b47ccad1c57c05912637e107096ba230c92b97187db79e19e},
  '{341, 1'b1, 512'he2fc500440f25769bdfcc82cca36025aa6e5335d8653935dee2cc2a8e8a37c8a886885663c7da8224d2e807f62e1f039ffffffff2aa58c5c932713706022af2a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h04452f554bae819b42effb84ef44a9f1cb7e2d75b4ba9ff9b9cfffaddde3fd1b, 256'h61a3fbc5e73c350f2e3d85a7452cd231a3f3375fc11f5fe153b185f53b09c1d0},
  '{342, 1'b1, 512'ha5ce1cdebbed43dea085a592a1ef6c0881660e99434c6f3d6ec24874bb6cc9d56400958f7f95fdc15d3dcc870056263b85ffffffff9f3ace8f83061d0410f802, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h05814f57f58efc7cb490119e584e635e6f0ad1c19fb5dc2edafda075bb55f98e, 256'h9dd5c6e39009d67d965903ecffe08a851775cc1248cc19c0b77798282131b8f6},
  '{343, 1'b1, 512'h6ea638f8043673b9b6a79ff39b5d311774de5f4d697e5251ede52feecabba85d705f25c58b7c2efc844ce598d1428d22e4b3ffffffffc75b0ecb7283d80278f0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdc1c4a46085e198843b1f01980cd5e4a1ff6f8e8ff7014397f0afd5b247fb0a0, 256'h38a13dc723ed90b30251d742b14733a03292ff26530a1ebcaf3d10862a6eff82},
  '{344, 1'b1, 512'h7cd22c5fec3646707603f858ccd785676b3284b63652913e5581a60e0c262034285489fb945534b7f2578b3e64e7b956bb6586ffffffffc05edada940cffb928, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1067667bf525734ca7f2510e36348fd9c2c9bccf032dfd571de6d45abd49361a, 256'hfa762568d3a19e5a1d8ea65e00202a5b16f9afae56733a01f86e35378c558da4},
  '{345, 1'b1, 512'hd289f68304c484efc5008425cbf00039a52c7b9d15476d36d58f1515d48a9ec94a850c121249365d7226fb6aad3a82c9eafe994affffffff58e8d36e4237022b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'he58d69dc56bc1031644847e3e046e2ea845a515d969d07ea1aa53aea5bd92fa1, 256'hbfe50b80f7c512f5ab521fe7e1a131045fde78d4de826c91573baaba1e35ca97},
  '{346, 1'b1, 512'h792eae16afd3069393b20db2ed2e192ffd845b08e10d076d8eafc98744329d6279d31d55ad56a090712fe131358feb130a94bc4a2fffffffff97daeec1130838, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hfe79c6b8c14d0f23d426e3d157f1b541f6bb91bf29957ef97c55949c9ba48a35, 256'h9da112c4a4cf4b1ff490c426f6c8ff122183964a0de56f7336ab382dc9d10285},
  '{347, 1'b1, 512'h51ae80a63d993770d8a5957111af53dabdf3abb9cf9908bc162ded716d3b3c5af2924c076e87c96249a4d7650253ff5112f8a2e7d2aaffffffff66e0e9175efa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h45d4ed7e9edacb5a730944ab0037fba0a136ed9d0d26b2f4d4058554f148fa6f, 256'hf136f15fd30cfe5e5548b3f4965c16a66a7c12904686abe12da777619212ae8c},
  '{348, 1'b1, 512'h100c883756f36d7c944d934c08932a99a1c2eb9892cc39a13a80b22aadc526ad755265f9ebbc8d0c1ccd31240299c71604332ff56592b7fffffffff1224308a3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4fb7c1727e40bae272f6143a50001b54b536f90233157896dbf845e263f24863, 256'h6fea5c924dca17519f6e502ef67efa08d39eb5cc3381266f0216864d2bd00a62},
  '{349, 1'b1, 512'hf4272253af2b51df321249280f3f3e62fb1e4a4a556f88bf3d5ae20ac5cc3e035e7b2141f9139b2f21d431068b8d5d96fcaad0f106289298ffffffff51777f01, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h779aac665dd988054b04f2e9d483ca79179b3372b58ca00fe43520f44fcb4c32, 256'hb4eca1182cd51f0abd3ea2268dcda49a807ad4116a583102047498aa863653f5},
  '{350, 1'b1, 512'h8bfa5531067a5cbc9bf002be2397bd10dd183d7ae47a02c0d0a7d87e1f94af93ea7365b711cfa611750ac963de0551c900dbad9cd8071b503afffffffffe6b6f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdb7ac6f65fb1c38d80064fd11861631237a09924b4eeca4e1569fa4b7d80ad24, 256'ha38d178d37e13e1afa07a9d03da025d594461938a62a6c6744f5c8f7d7b7bb81},
  '{351, 1'b1, 512'h8a5409853b325b917b8a2aa1eb394767bb07fa82af11357e777f7404e0955bc9bb9cc5a918475c52df4772a1207e3ee4f3e3d3c8e68e84e10477ffffffffd35f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hc90043b4aadf795d870ac223f33acdbd1948c31afff059054dc99528c6503fa6, 256'h829f67b312bb134f6954a23c611a7f7b5b2a69efced9c48db589ac0b4d3da827},
  '{352, 1'b1, 512'h8e38a571ec826b9af00de0c523b6e073aaf9380cc64fbc86755f33f065361d8963ea2c42796ac7516f53d689e1da364bb7caf6b22a5fee81410646ffffffff7f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hfa16c0125b6615b90e81f7499804308a90179bf3fcff6a4b2695271c68b23ded, 256'h0d6cda5ce041dc5a5f319ad9c0de4927d0cf5e89e37b79216194413d42976d54},
  '{353, 1'b1, 512'h0f3ad12803aaf9bc615745a47da85dd90bff191d3e9441cc2cc96bf8c01f5e514b256685e3e48f01a98a5f27d20cd1c317a6f816ca8611fbc8891236ffffffff, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1a4b5bd0f806549f46a3e71bfe412d6d89206017640ded66f3d0b2d9b26bec45, 256'haac5f74e3130264e01428570ee82ee47e245d160ed812ae252dedffd82e1ec2c},
  '{354, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 256'hc7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hf8e272234b51475ec4c6f327562a6e5c9080a96225e88b2e5f72a8eecbd41ab4, 256'h516b91617fc39e3141b3bc769f6a3b2e468e687f50bdc29e19088af62d203f4b},
  '{355, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hb6e08b1bcc89e7fb0b84d7497e310553495be4877eccc4b3d6d79f7c68a05734, 256'h31760fa1bcea4972759174ac1103bc6011985ccee251918d0573fbcb78969116, 256'h000000000000000000000000000000004319055358e8617b0c46353d039cdaab, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},
  '{356, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hb6e08b1bcc89e7fb0b84d7497e310553495be4877eccc4b3d6d79f7c68a05734, 256'h31760fa1bcea4972759174ac1103bc6011985ccee251918d0573fbcb78969116, 256'hffffffff00000001000000000000000000000000fffffffffffffffffffffffc, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},
  '{357, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h3590c6a10353d669bc94d8e2ff9e14bbeed4a7f45b887255ab7e37b676387bb6, 256'h15fc6f97ce39a3874c2b34cc571889abfa0a706c2cfb0e5a4750cc25690696f8, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254f, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},
  '{358, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h369e96402f2cfd1a37b3acbdecfc562862dbca944a0f12d7aaacb8d325d7650a, 256'ha723621922be2bdac9186290fdcdda028d94437966507d93f2fc1f5c887fdedb, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h909135bdb6799286170f5ead2de4f6511453fe50914f3df2de54a36383df8dd4},
  '{359, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h27a0a80ea2e1aa798ea9bcc3aedbf01ab78e49c9ec2ad0e08a0429a0e1db4d0d, 256'h32a8ee7bee9d0a40014e484f34a92bd6f33fe63624ea9579657441ac79666e7f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h27b4577ca009376f71303fd5dd227dcef5deb773ad5f5a84360644669ca249a5},
  '{360, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h9cff61712d4bc5b3638341e6e0a576a8098c9c6d3f198d389c4669f398dc0867, 256'hf3b9e09f567f3dfd9c4d2c1163e82beadf16c76e8f9d7a64673800ea76fa1e59, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{361, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hd9117cae81295e82682fa387991e668e1570e0e90100bf4e63964822460561bc, 256'h19f96b1787ed15769929978ba3dd7f68c97adf5c16f671e756cd8f08c49456ca, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000003},
  '{362, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h8cfcbad3524c22b992529f943e3ce0b2d126085501d6e3edd4f1dbf74bdca21e, 256'hafb259b1ba179cac09e8e43a88c8a09e7339910a7c941932e44b8be56f1fccde, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000005},
  '{363, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hfbb51127e1f1b6a38e9fe9a2544614edb8e43ad7cd8c56f14b3235dda3bc1117, 256'h9abd9753a9e647e9340c395fb2b91384d6d33fcb6456214350b6f3fa00f4364c, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'h0000000000000000000000000000000000000000000000000000000000000006},
  '{364, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hfbb51127e1f1b6a38e9fe9a2544614edb8e43ad7cd8c56f14b3235dda3bc1117, 256'h9abd9753a9e647e9340c395fb2b91384d6d33fcb6456214350b6f3fa00f4364c, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632556, 256'h0000000000000000000000000000000000000000000000000000000000000006},
  '{365, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hdc80905500d7d74ed47de5224d8734545f22b776ae086cabfffe6ce58d5ef994, 256'hdc3067ce7d2cdfa9f4d5ace296b752814acc69c19a932d8b14077927901de3bf, 256'h0000000000000000000000000000000000000000000000000000000000000005, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc75fbd8},
  '{366, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1b824a11eed94fbcd9b722d06613bbcf7eca00b9136f2652642178f37b1a920e, 256'he900de495d9ef56fa6d19f3dd1e0edb23d23835ac8c2d3d13c0227e852e503eb, 256'h0000000000000000000000000000000000000000000000000000000000000100, 256'h8f1e3c7862c58b16bb76eddbb76eddbb516af4f63f2d74d76e0d28c9bb75ea88},
  '{367, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2914b30c4c784696ffc3dddcec05f36cb1488bc342b9f529d5387acb9e48cb8d, 256'h3dbd30d0d5d6d6a39108863c2d6a6e8571cd3261fb9eb98ce46125bd8f139136, 256'h000000000000000000000000000000000000000000000000002d9b4d347952d6, 256'hef3043e7329581dbb3974497710ab11505ee1c87ff907beebadd195a0ffe6d7a},
  '{368, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2579f546fe2f2aeb5f822feb28f2f8371618d04815455a7e903c10024a17da41, 256'h5528e951147f76bee1314e65a49c6ec70686e62d38fbc23472f96e3d3b33fd1f, 256'h000000000000000000000000000000000000001033e67e37b32b445580bf4eff, 256'h8b748b74000000008b748b748b748b7466e769ad4a16d3dcd87129b8e91d1b4d},
  '{369, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hb102196bf455ee5aafc6f895504d3c3b6b2d37c35f8669bd0f0b694795fbd992, 256'hf777b6f829b9628ac35db0ef43f6a89f0a42812614e4c15924d8d47ebe45bae5, 256'h0000000000000000000000000000000000000000000000000000000000000100, 256'hef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},
  '{370, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4d056ab2ff57662fd6eebbe23930fef5cd08083e24146190cd01960b1fcd3749, 256'hfe7ec5847651c857898be0f09efd6e0116a5dbe327f6f3080a65fc966bf64d91, 256'h00000000000000000000000000000000000000062522bbd3ecbe7c39e93e7c25, 256'hef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},
  '{371, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h361c4a62cd867613138dfe24ccebc4b7df1b55fc7410f4995ee2b6b9ab222058, 256'h4f116c6c84e53d262fd13a5f5de6b57e7a1981de4ecdffdf3323b4e91d80649c, 256'hffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc6324d5, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},
  '{372, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hdb9d5c5113f00822a146c9cda2e75cb6634cd0dff54aff6e22875171f57a0dad, 256'h1c424cdd83eb01c02f6f8d36f42c6dc7e39db74358da8ac9bc9dc5890d46f667, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h0000000000000000000000000000000000000000000000000000000000000001},
  '{373, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hdb9d5c5113f00822a146c9cda2e75cb6634cd0dff54aff6e22875171f57a0dad, 256'h1c424cdd83eb01c02f6f8d36f42c6dc7e39db74358da8ac9bc9dc5890d46f667, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{374, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h99f19f07b33e03caf4703e04b930d57d6d9baa44460c596a2d3064e0b63ea412, 256'h86a74c4612a812ee348d2b43f80de627c11c75d81511e22a199c32119b792c6a, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},
  '{375, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h313f3309b236484c6eb4ea381e007854467a617343a2e97d845801c01a632cfe, 256'h33f231854bba89a8ca3f802a2764d3bf6c3233c811a31e5e8028a0b862cb1977, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8},
  '{376, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hd3aa01fe59bad92cffe3db59e1385391fafd7af4e4ce462e8aac157274cc8a05, 256'hc7a7e603e18538aac15f89610beacc21e39898e6c5f7680a81c5bd7bd744a989, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9},
  '{377, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h5e31eccd4704ebf7a4247ea57f9351abadff63679f2276e2a3b05009ebc1b8df, 256'h648465a925010db823b2a5f3a6072343a6cc9961a9c482399d0d82051c2e3232, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281},
  '{378, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hce0a47f881fd7315a733c4317848fa33c72e38de0b8fda36b61aa9a164f5808a, 256'h85b05d25115ea4097ddf63f878c8e83657e66de136a8f9e62ed81a58bf117ff9, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'hbc07ff031506dc74a75086a43252fb43731975a16dca6b025e867412d94222d0},
  '{379, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hcd6f487b47f36c0dea8f4b04c4e6ac637c76b725929c611f48addcf3d2f65941, 256'hb50ea8f3a491190ee0b20cfb6efd113608e7c7c127577500e7f5c4a4e490fd60, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},
  '{380, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h456e5f8067d68a1b0a2e8fe2b28acad5755687154a0f167734ebabbdc059070d, 256'h720dbe96659a66ef0cf27a73e7b3f3f145a60e0ad29f1e21dcc2bb42f0d82c1e, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'haaaaaaaa00000000aaaaaaaaaaaaaaaa7def51c91a0fbf034d26872ca84218e1},
  '{381, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h42bf0c0ac1e3850baf5515748a878e34249f71035e20a9f54ed468ec273cb0fc, 256'h5b3138500230055c71f12d53f5c7d0e3d8aa54a94c668cb311e20d195fc71abb, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h6bfd55a8f8fdb68472e52873ef39ac3eace6d53df576f0ad2da4607bb52c0d46},
  '{382, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hffdd48da63d3af67223f16c51eb7e95600eb0b0e8b964f4fcd8c534face3c2c2, 256'hb4e009ab2a76829480e69c9e43b2f1fe076cfafb3fa8d27dd4d6bab4d6c3db54, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h654937791db0686f712ff9b453eeadb0026c9b058bba49199ca3e8fac03c094f},
  '{383, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h793cbfce6f335dcfede7c6898ea1c537d7661ed6a8c9d308d64a2560d21c6e2c, 256'h483d23a5ff05da00eaf9d52cf5362be9b53b95316c6a32e9ebe68d9ac35c2fd6, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hc51bbee23a95437abe5c978f8fe596a31c858ac8d55be9786aa5d36a5ac74e97},
  '{384, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'ha9f7023f559d4bb6c9f4bc3643e2824aff5451d929479ec3ea5eb30bad2c36ac, 256'h6a7c77e8dd21f4ad49b103e67da9d3cda62b653dd194fad2ba8d1dd37bb0ea9b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h8ba4c3da7154ba564ab344ae12005aa482b6c1639ea191f8568afb6e47163c45},
  '{385, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hdf79ee082b2fc77e9ce4633471f569bbcb5ce53856e3067774f37e8a64a2c7ff, 256'haa488a6c34d499df76f427de3609bfcfd9feae67ffe0b0de594463c453b0ab16, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h4c3dafcf4ba55bf1344ae12005aa4a74f46eaa85f5023131cc637ae2ea90ab26},
  '{386, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4cc3bf65e32e00284adfca00f40df755415c485091ac0489ae9a337103a5f8f0, 256'h123ab86dd433b933b4f2063c002144df3cfeba78dad0ed89c0377541532908c2, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h987b5f9e974ab7e26895c2400b5494e9e8dd550bea04626398c6f5c5d521564c},
  '{387, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h264a7ad439a4828a9dc97ecf837155355f99ae0b65975f851b541ad3a0e032f0, 256'h67268b7298c73e581866fbcbd161689b16b81cf262e007ce68e25a28c83ef041, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hfcf97e2fbf0e80d412005aa4a75086a3f004f59d512cb47271798733ab418606},
  '{388, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1d7ff4d3a41206c8143635f12876e0ea0875ea5e4a5a249250d0eda33daa211f, 256'h56e89c0beaf910ac934ca12380455600d0fd85b56a7035cb171b3f1c72a15569, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h79d482b60864d6c5cb4fd5db9e7e28ccd9a5948c316c8740fb429c0f37169a02},
  '{389, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hb09685f338dceb421778a1458d52bed734c236242da2baa280d6f6b7b86e4f11, 256'h7fe6a34146b422d7aebd1a51b20948d7872a514c4cfd7686dc436b70733d6473, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h8ecd11081a4d0759c14f7bf46813d52cc6738115321be0a4da78a3356bb71510},
  '{390, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hdd811f2c0f5e9d4fbb2ef31818c1cd807247bc14fcd1170bef00e2c71dc037b4, 256'h43a15cdf8f3fbdc87e06250c0720d261d2b8d087fa7bf9548f6293f0ce5ae899, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'he8dbffed13c9a2093085c079714f11f24eb583d73ba2b416b3169183e7d9b4c2},
  '{391, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h69d60ae1f39e1da95809d408894707ad2134f4943a1db089bebf815a391f18db, 256'h32b401d98bf894d3b6d59e6eb45573285642e358ad687b7d7bf9600b1987809e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hca01552a838124bec68d6bc6086329e06673900eac5c262e5ce79a8521cd1eae},
  '{392, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'ha658553a0620c95e987b5c3163bcfea68c52065f53c9d553f2a924d8b3ed511f, 256'h79f0dfec4536b65aa5fb31297e96f6b464aa669b9268b3156c43d4612978a577, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h9402aa560702497c8d1ad78c10c653c11000256fb1a0add7c6156a474737180b},
  '{393, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hbc4d3354a6a973dd8088919cc181194e879ed7920db30d0d1278edf74413b7b9, 256'h2450d162b26dcb25fbbd53ea4044189981d737055925bd2e86bfb0374b09f3ca, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5e03ff818a836e3a53a8435219297da1b98cbad0b6e535812f433a096ca11168},
  '{394, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h0eb628724fce764c687d874ade7b8e0aa4abf20ee6e3610fac9fe3e72f97ab5a, 256'hed09f4843660eb1daf015d397a7c1073d7ae43bda0ba3e117008785abfffa00f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'he28ddf709d4aa1bddf2e4bc7c7f2cb516cb642bb3e39c3feaf2fcf16ab9539f4},
  '{395, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'he7ac5cc7f296912f703f59fe88e49b521da245e12e6eee161ee6b3b1127611a7, 256'h7b3bedd2a773cf58b0629b936dd85dad2d0c39676306ed63e1a9bcd0e08bccc2, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffffaaaaaaaaffffffffffffffffe9a2538f37b28a2c513dee40fecbb71a},
  '{396, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2407b60abf3ee5edaf92ed505a11d0ddce0ea33eca58a031bb2f162c512f4062, 256'hfb81bff36bf967e834e3d5d468730dcd70440022ab60061a62fac53350fe259f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hb62f26b5f2a2b26f6de86d42ad8a13da3ab3cccd0459b201de009e526adf21f2},
  '{397, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h47b2ad96dfc2f23fe5926809f38042b2c801962bd7394cefbf4aacb2554b7b0b, 256'hdf2b937a16a7d96a2a0682cd164428890208597f2cdcc734fda73600b5cf6c59, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbb1d9ac949dd748cd02bbbe749bd351cd57b38bb61403d700686aa7b4c90851e},
  '{398, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h69a65b75f31ae7b4930292f90902461befcee5d1606939c28e01b652a7fbc498, 256'hcf68619e5860128f56cecf53eba2ffe82889a9bb04a5fa4c8b722bc91d55978a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h66755a00638cdaec1c732513ca0234ece52545dac11f816e818f725b4f60aaf2},
  '{399, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hb2037176c84db04a6c773e32f9ed1d6b25ef4c303c6725c6932ec2cc2788bcbb, 256'h9361505e6b771691adb41598f292d6521722404bf183241b195738b77abd6cfe, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h55a00c9fcdaebb6032513ca0234ecfffe98ebe492fdf02e48ca48e982beb3669},
  '{400, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1eef95aef71f793afd50bb2604064d63e88bef7404a4d0e206446245ae2e7834, 256'hc96e86dd040f9794b63712d90e719576b8b92c406ab0f288ad9b327bd124454f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hab40193f9b5d76c064a27940469d9fffd31d7c925fbe05c919491d3057d66cd2},
  '{401, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'ha9734899c954e5b7adbca8f783428b5fbcbdfd3d2813f8d2f95b31a78ab10756, 256'h7667abf8c02ce4951bc59b2564130c27d7b64cdbc5cad95ca42d5bbb7cd4e793, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hca0234ebb5fdcb13ca0234ecffffffffcb0dadbbc7f549f8a26b4408d0dc8600},
  '{402, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1ae51662331a1dbfab0751d30dfab2273a04a239e055a537b16ab595f9612396, 256'h434f21c2bfe6555c9fc4a8e82dab1fa5631881b016e0831d9e1bbf5799fcf32e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbfffffff3ea3677e082b9310572620ae19933a9e65b285598711c77298815ad3},
  '{403, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h53c90cdd8b0dadd21c44ad557b327f4dbf57144aaf06597deb3f94125206a6c1, 256'h4603475bd79b30e36340cd09b0b59e6cd46ce90150e9ffe5c8a0172b2c9898e3, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h266666663bbbbbbbe6666666666666665b37902e023fab7c8f055d86e5cc41f4},
  '{404, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h33797539515c51f429967b8e36930d9fdda1edb13aecec9771f7cde5f6f2e74e, 256'hba51d0b6456bb902dba1f3ea436f96ad2355da454dc9b32c503c4bc6cfd6d410, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbfffffff36db6db7a492492492492492146c573f4c6dfc8d08a443e258970b09},
  '{405, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h0a8f5f1d5bbd2783fa7f37c86879057fb2fcf25383aafb86d03d6bafb41a17b3, 256'heaf6da715fe950349fd5736117b08e15e32cf1d2fdc003e510009f1b4ba1e648, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'hbfffffff2aaaaaab7fffffffffffffffc815d0e60b3e596ecb1ad3a27cfd49c4},
  '{406, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1dbc94e96c056b9d2cb6773bb24b69ed473851badf927a29955aff290ef3675a, 256'h65e587561122aa8226facb95df08308cadf01c8351a1569176d917821113aa7c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffff55555555ffffffffffffffffd344a71e6f651458a27bdc81fd976e37},
  '{407, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h084ab885dbff7f12e6cdadb59d456e500797779425c7518c259c83718289e6e9, 256'h91c345d3a093e86670605bbc2ff4c69d0ed694fd433ec6b6ba1bf7d56c3e6b51, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h3fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192aa},
  '{408, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h003adfa4c620a207096cd18ee8fd2a90e20106cf824a0c63d6dec727a9fe7f50, 256'h9430d26bdd5f71e819d12b70069901461ae083cc809122d4fb86b5c475244e5a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5d8ecd64a4eeba466815ddf3a4de9a8e6abd9c5db0a01eb80343553da648428f},
  '{409, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h7c98b2d47eb433c0d18e533cfbc8909d66f7b79d5925ccb17eccec9d105c5884, 256'h8d5ca99b350bd7d10ab5ee6fcfe46623fdc03e9f828158f4d4cc08ad1ff83de4, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 256'hb4cfa1996ec1d24cdbc8fa17fcabc3a5d4b2b36cf4b50a7b775ab78785710746},
  '{410, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h7c98b2d47eb433c0d18e533cfbc8909d66f7b79d5925ccb17eccec9d105c5884, 256'h72a35663caf4282ff54a1190301b99dc023fc1617d7ea70b2b33f752e007c21b, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 256'hb4cfa1996ec1d24cdbc8fa17fcabc3a5d4b2b36cf4b50a7b775ab78785710746},
  '{411, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hb7a90e21e7547d73267940033cea05042c50f7c9fa5eaeb471cd6260c685f2e3, 256'h8bb7309d0c3bab249faaf3e44179d6dd5302375c580fd0570a788c6be3680c67, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},
  '{412, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1550a173373b2d594374f0642cd73de06a045c09c7a4f388c731e8cd8971adfc, 256'h9a3a9843583a86c0e1c62cbde67165f40a926b1028ba38aa3895e188ebbc7066, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // OUT_OF_RANGE r_len=33 s_len=32
  '{413, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h313447778195daa1791a6530cd0697ae34bf9d8d225984394f72eef350597111, 256'h0996a8fbdd1a70ecd64cb00b595afe1669bfef80d91756a62d84c1d83e0f22ab, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},
  '{414, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4ada634941476ca63c2c5803eec2f33b2d17920f798a5be6275f5a54cd2e7639, 256'hb1a04bead5c7314c427492db21b9544d81caa8159587e41aa023aa967f31aaa1, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},
  '{415, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'haacce093270fa59ad412b5459a08e490743b97086c781ac3c8d54030b41a3119, 256'h3bece4956172d56befb7011d684e772905e48d2115444a75ac7a325a3f25f4b1, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'hb6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},
  '{416, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hf62b8d7feeff5a847ab79212269e55e62fa87ebe930821747b57a511a5ea99f0, 256'h439ee057bb27898582a683c3fdb7f95404d41d42f276803751a316eb3aab7ebf, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'hcccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},
  '{417, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4baa07ff6e7bb9aa223d1c61932005fe98fe78b787fdab4bd3619bc8833072a2, 256'hbcacd63802c56af82607953e72a0f5d3c23bd265544e020951824ea485555d33, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},
  '{418, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h0c753ed1ba92f766800fdd0ae1c0d7f8f4cd8305fd803d8bca881397b5937e2d, 256'hb568509b1faf3cf251de6db9810e8b8caed235da10eeddbed62775c8e5c9460a, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},
  '{419, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h030fdcae6541f22c5bab254e4f1a285c507d1cefea03bf90cf19daf3cb62df69, 256'h5ff2c94d588f2c2b2b0a12bebc011bcee4fa1b54506ec07d0a29d24a0891193c, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},
  '{420, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h03fc621eaf90c23d8f9fa125d2c59b8728ebccb30ca3e3db879a06ca90f20cdc, 256'hae58d3f0c6aef0e805be10ea54e23cf6f0397f9addddc2b09088855316b0ef44, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},
  '{421, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h70f2ce24dc62923bb09cc92d74329bbd0d2e6b0e354c0be2383d24acdccb9e4c, 256'hd42d1f973466f5e5462a939084a294ebfc7a45629c70ee5def46de9536ea7bf7, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'hb6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},
  '{422, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h732b8ac0c30fe44307431235271cb5d6e5f677a19ce3f058b939a7bf19349d3c, 256'h858cc735af8577468275847cf5ec19972e6c20738276e2708b23c595bfc4433d, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'hcccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},
  '{423, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h47aff9501825a166782bb58a5b459006eacdbce5e5323addad34ec1b6444cdce, 256'h9199c31502ad4277c73ddd0c807b72634c45762404837d9814a5d4b5a7c3f398, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},
  '{424, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'haed8eeff77644bf83b9222f8f57173fa8217ec7e0763ee7d7171fb6092fba5c0, 256'h6486a86d94f48834ba5adbaf349687f9cee400389642b828e68207b147ca2c46, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},
  '{425, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'hf7c54a585a904300d05b53ef3b854e71999a344b89adc0caaa28e254db9bc7c7, 256'hc161a79f38ff446051303577e40638fb020329940a63c241bb32c2205eb57b7d, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},
  '{426, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},
  '{427, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'hbc07ff031506dc74a75086a43252fb43731975a16dca6b025e867412d94222d0, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},
  '{428, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'hb01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},
  '{429, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'hb01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'hbc07ff031506dc74a75086a43252fb43731975a16dca6b025e867412d94222d0, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},
  '{430, 1'b1, 512'hcf83e1357eefb8bdf1542850d66d8007d620e4050b5715dc83f4a921d36ce9ce47d0d13c5d85f2b0ff8318d2877eec2f63b931bd47417a81a538327af927da3e, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 256'h87d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h093f3825c0cf820cced816a3a67446c85606a6d529e43857643fccc11e1f705f, 256'h769782888c63058630f97a5891c8700e82979e4f233586bfc5042fa73cb70a4e},
  '{431, 1'b1, 512'hdc5e71048a56da7aa1bf5fad1ae227446663488d8a531d490c4b5efa048ca4651acd9a196d9b13ee2a1c74ad440bdd88f6a34a02fbfadac2f7ce869e64486558, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 256'h87d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'he8564e3e515a09f9f35258442b99e162d27e10975fcb7963d3c26319dc093f84, 256'hc3af01ed0fd0148749ca323364846c862fc6f4beb682b7ead3b2d89b9da8bad4},
  '{432, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 256'h87d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h1412254f8c1dd2742a00ddee5192e7baa288741026871f3057ad9f983b5ab114, 256'hbcdf878fa156f37040922698ad6fb6928601ddc26c40448ea660e67c25eda090},
  '{433, 1'b1, 512'hd296b892b3a7964bd0cc882fc7c0be948b6bbd8eb1eff8c13942fcaabf1f38772dd56ba4d8ecd0b626ff5cef1cd045a1b0a76910396f3c7430b215a85950e9c3, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 256'h87d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h9e0676048381839bb0a4703a0ae38facfe1e2c61bd25950c896aa975cd6ec869, 256'h6ea0cedf96f11fff0e746941183492f4d17272c92449afd20e34041a6894ee82},
  '{434, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 256'hed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h554482404173a5582884b0d168a32ef8033d7eb780936c390e8eedf720c7f564, 256'h0a15413f9ed0d454b92ab901119e7251a4d444ba1421ba639fa57e0d8cf6b313},
  '{435, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 256'hed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h0b1d838dd54a462745e2c8d5f32637f26fb16dde20a385e45f8a20a8a1f8370e, 256'hae855e0a10ef087075fda0ed84e2bc5786a681172ea9834e53351316df332bbd},
  '{436, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 256'hed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'haf89e4f2b03e5d1f0352e258ef71493040c17d70c36cfd044128302df2ed5e4a, 256'h420f04148c3e6f06561bd448362d6c6fa3f9aeeb7e42843b4674e7ddfd0ba901},
  '{437, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h84fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h6c1581f1485ccc4e657606fa1a38cf227e3870dc9f41e26b84e28483635e321b, 256'h1b3e3c22af23e919b30330f8710f6ef3760c0e2237a9a9f5cf30a1d9f5bbd464},
  '{438, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h84fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'hdc83bf97ca28db0e04104a16fe3de694311a6cd9f230a300504ae71d8ec755b1, 256'h64a83af0ab3e6037003a1f4240dffd8a342afdee50604ed1afa416fd009e4668},
  '{439, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h84fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h575b70b4375684291b95d81e3c820ed9bde9e5b7343036e4951f3c46894a6d9d, 256'hf10d716efbfeba953701b603fc9ef6ff6e47edef38c9eeef2d55e6486bc4d6e6},
  '{440, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h8d4f113189dfd3d3239e331f76d3fca9cef86fcd5dc9b4ab2ca38aeba56c178b, 256'h78389c3cf11dcff6d6c7f5efd277d480060691144b568a6f090c8902557bfc61},
  '{441, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h834d10ec2d2d50eeebfecd6328f03fafbb488fc043c362cbc67880ec0ebd04b3, 256'h94c026feaf6e68759146fe5b6fd52eaa3c3c5552d83719d2cb900615e2a634db},
  '{442, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h6894de495e7bb5566807d475d96a0d414a94f4f02c3ab7c2edc2916deafc1e1f, 256'ha603642c20fabc07182867fcc6923d35be23ad3f97a5f93c6ec5b9cce8239569},
  '{443, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 256'ha01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'he500c086fedd59e090ce7bfb615751ed9abe4c09b839ee8f05320245b9796f3e, 256'h807b1d0638c86ef6113fff0d63497800e1b848b5a303a54c748e45ca8f35d7d7},
  '{444, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 256'ha01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'hb922c1abe1a8309c0acf90e586c6de8c33e37057673390a97ff098f71680b32b, 256'hf86d92b051b7923d82555c205e21b54eab869766c716209648c3e6cc2629057d},
  '{445, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 256'ha01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'h823c37e46c74ec8497d89245fde3bf53ddb462c00d840e983dcb1b72bbf8bf27, 256'hc4552f2425d14f0f0fa988778403d60a58962e7c548715af83b2edabbb24a49f},
  '{446, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hfffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h577a08a95db6dcda9985109942d3786630f640190f920b95bd4d5d84e0f163ef, 256'hd762286e92925973fd38b67ef944a99c0ec5b499b7175cbb4369e053c1fcbb10},
  '{447, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hfffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h7ba458cfe952326922c7aa2854bdc673ce3daaf65d464dfb9f700701503056b1, 256'h0df8821c92d20546fa741fb426bf56728a53182691964225c9b380b56b22ee6d},
  '{448, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hfffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h5cd60c3b021b4be116f06f1d447f65e458329a8bbae1d9b5977d18cf56184861, 256'h4c635cd7aa9aebb5716d5ae09e57f8c481a741a029b40f71ec47344ef883e86e},
  '{449, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h00000003fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h4b50e1e8cf830e04c17e7472caf60da8150ffa568e2c64498cc972a379e542e5, 256'h2e3adaa5afab89cca91693609555f40543578852cde29c21cb037c0c0b78478e},
  '{450, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h00000003fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h5aea930c7d8fffcd5c6df2c9430ef76f8b5ed58a8b9c95847288abf8f09a1ac2, 256'h7ddfef7688a6053ce4eeeeefd6f1a9d71381b7548925f6682aa0a9d05cf5a3a3},
  '{451, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h00000003fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h98b092c2d14b5b14a23e9368e0ce1be744dfae9f9a5cdaba51e7872099df96f2, 256'h90d3e4f87bd7bc94589f8150b6b01045cd8759a00af78b24d7de771887610df5},
  '{452, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hbcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 256'h000000001352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h9e95f2856a9fff9a172b07817c8c60fe185cd3ce9582678f8cc4b02bc444621a, 256'hc54ca51d8117d904f0d3773911cb2792348fae21c2da7dad25f990d122376e4c},
  '{453, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hbcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 256'h000000001352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'he77df8f9782696344c33de29ebdc9f8d3fcf463d950cdbe256fd4fc2fd44877e, 256'h87028850c962cf2fb450ffe6b983981e499dc498fbd654fa454c9e07c8cb5ca8},
  '{454, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hbcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 256'h000000001352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'hbd2dd6f5026d2b5ad7ead74bdf52b8cbcabc08facee0a1c8584658a85ed0c5dc, 256'h3e8543e819bdae47d872e29a85ba38addf3eaeaad8786d79c3fb027f6f1ff4bf},
  '{455, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hbcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 256'hfffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'hbd5c0294acc28c15c5d1ebc7274c9ca21a081c8a67da430a34a7fff1a564fabb, 256'h7ec103a2385b4ff38b47d306434e9091de24dc9f1a25967ee06f8a0a53ac0181},
  '{456, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hbcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 256'hfffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h3c7dbfb43dd80379ee2c23ad5472873a22c8a0179ac8f381ad9e0f193231dc1f, 256'h7cf8e07530ade503b3d43a84b75a2a76fc40763daed4e9734e745c58c9ae72d3},
  '{457, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'hbcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 256'hfffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'hb38ca4dac6d949be5e5f969860269f0eedff2eb92f45bfc02470300cc96dd526, 256'h1c7b22992bb13749cc0c5bc25330a17446e40db734203f9035172725fc70f863}
};
localparam int test_vectors_secp256r1_sha512_NUM = $size(test_vectors_secp256r1_sha512);
`endif // WYCHERPROOF_SECP256R1_SHA512_SV
