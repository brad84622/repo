`ifdef WYCHERPROOF_SECP384R1_SHA3512_SV
`define WYCHERPROOF_SECP384R1_SHA3512_SV
typedef struct packed {
  int           tc_id;
  logic         valid;  // 1: expected pass; 0: expected fail (zero/oversized)
  logic [511:0]  hash;
  logic [383:0] x;
  logic [383:0] y;
  logic [383:0] r;
  logic [383:0] s;
} ecdsa_vector_secp384r1_sha3512;

ecdsa_vector_secp384r1_sha3512 test_vectors_secp384r1_sha3512 [] = '{
  '{1, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'h302d08b563b09fbd4bb648f56a35794a12d24f48cefb874eac860c115c043020c92da2a8a55ad7b52aa165bbb90ff909},
  '{2, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{3, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{4, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{94, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab760000, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=50 s_len=48
  '{95, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hf74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a0000},  // OUT_OF_RANGE r_len=48 s_len=50
  '{99, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab760500, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=50 s_len=48
  '{100, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hf74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a0500},  // OUT_OF_RANGE r_len=48 s_len=50
  '{115, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // r=0
  '{116, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{119, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=49 s_len=48
  '{120, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=48 s_len=49
  '{121, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7abf6, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{122, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b530ea},
  '{123, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h00fbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{124, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'h00cfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b530},
  '{125, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=50 s_len=48
  '{126, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=48 s_len=50
  '{129, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // r=0
  '{130, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{131, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e0318ffb708876bbed3734ce2578a5d7d5a7c049163f7cd4e9, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=49 s_len=48
  '{132, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e0a2c9606ca008602e8700b2c0e74488dfcde81640a5f28203, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{133, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h042dc5e4fb2d96936337926c3717cdabd87fd0188ef09a1f95d352116bc071f220e53f8cd00acfa5452bd0548d48548a, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=49 s_len=48
  '{134, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h042dc5e4fb2d96936337926c3717cdabd87fd0188ef09a1f5d369f935ff79fd178ff4d3f18bb77203217e9bf5a0d7dfd, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{135, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h042dc5e4fb2d96936337926c3717cdabd87fd0188ef09a1fce70048f77894412c8cb31da875a282a583fb6e9c0832b17, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=49 s_len=48
  '{136, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=49 s_len=48
  '{137, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h042dc5e4fb2d96936337926c3717cdabd87fd0188ef09a1f95d352116bc071f220e53f8cd00acfa5452bd0548d48548a, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},
  '{138, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b0e2408ef28c6a2b9de70678bbec067740af36cd19e07a59dd},  // OUT_OF_RANGE r_len=48 s_len=49
  '{139, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b15379f3eea3fbcfdf36d25d575aa5284ad55e9a4446f006f7},
  '{140, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'h302d08b563b09fbd4bb648f56a35794a12d24f48cefb874ee522be8f67cd0241711394f65caa303a3db54c50ec4acf96},  // OUT_OF_RANGE r_len=48 s_len=49
  '{141, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'h302d08b563b09fbd4bb648f56a35794a12d24f48cefb874f1dbf710d7395d46218f9874413f988bf50c932e61f85a623},  // OUT_OF_RANGE r_len=48 s_len=49
  '{142, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'hcfd2f74a9c4f6042b449b70a95ca86b5ed2db0b7310478b11add41709832fdbe8eec6b09a355cfc5c24ab3af13b5306a},  // OUT_OF_RANGE r_len=48 s_len=49
  '{143, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbd23a1b04d2696c9cc86d93c8e8325427802fe7710f65e06a2cadee943f8e0ddf1ac0732ff5305abad42fab72b7ab76, 384'h302d08b563b09fbd4bb648f56a35794a12d24f48cefb874ee522be8f67cd0241711394f65caa303a3db54c50ec4acf96},
  '{144, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // r=0, s=0
  '{145, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},  // r=0
  '{146, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},  // r=0
  '{147, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},  // r=0
  '{148, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},  // r=0
  '{149, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},  // r=0
  '{150, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},  // r=0
  '{151, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},  // r=0
  '{154, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{155, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{156, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{157, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{158, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{159, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{160, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{161, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{164, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{165, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{166, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{167, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{168, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{169, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{170, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{171, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{174, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{175, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{176, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{177, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{178, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{179, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{180, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{181, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{184, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{185, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{186, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{187, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{188, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{189, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{190, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{191, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{194, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{195, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{196, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{197, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{198, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{199, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{200, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{201, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{204, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{205, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{206, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{207, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{208, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{209, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{210, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{211, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{214, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{215, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{216, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ff},
  '{217, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52973},
  '{218, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972},
  '{219, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52974},
  '{220, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000ffffffff},
  '{221, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff000000000000000100000000},
  '{230, 1'b1, 512'hb59b66a376f7e41f12114cc5359cb352c1390ce74c9e76a02ee4e1ebc58af0a2801b014036f29a20848a952718749f92efe909acec366c9e3c308614a4506d3a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hac042e13ab83394692019170707bc21dd3d7b8d233d11b651757085bdd5767eabbb85322984f14437335de0cdf565684, 384'he0f133f6ff3dd2496a15abc92b34315a17f49679734720c0270f5dad3dcd2833f913b48a6cdf2ec6b2ffc9d3d72d545b},
  '{231, 1'b1, 512'h0000000097ae34ada66084471ced074cb11f6012595501e4f88b5ab4526808fbaabfff3975c6cf53455cee950965a5b5b71310c8a1822cb5d15b513b43dc5720, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h202858607c9a8777f7001f0fb25b12f39d5fb1b86b767adb1a32fd8ca18dec71d0cf69a3839f3097d9132247b558e1b6, 384'hd7be6ca34d3a846195b67e5bb517fb169ed4da4ee124b854637c7f86bcacbad64caa4e9e50fb932c1679b463ffa87b23},
  '{232, 1'b1, 512'h4a00000000d34b9c928306129f1a8059b199049f30ffd4d5b9747c848b197497634fb5190298af2f6a90d273164d68431c984e0fcd3a810ccd7b95b5e0dcd21f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hbbd2e99974a733000592ebad069c39adcb4ee32718f262dc167fa0b4080e788c95cf177bcff61b72dcdf7406906af995, 384'h89552e369143d56a006b90b8b3fd68cdb49a8f26ec5ca4df03abc149273de0a4693af37362f3c689a6d8b6935663273e},
  '{233, 1'b1, 512'hf25200000000600b35bfa47958845baa9428119e3a1641db59a3b72db0b47470dc44921ca1826d81bc2e78142986441cb6a6c15880383e1ed77282f966ad17de, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb35e96f93302bc08e339bfbb2fbe04872f1eca413084629041ffc0dd94eee677bc32cb09022ed6214153f2ed705edb22, 384'h5aee1acff79c6bdbbb4d3c656c3010eba72fa671df68637a5fbbc2dd2268bbb4fef4a85c90b49013e0c1a2aecd342b6c},
  '{234, 1'b1, 512'h9e93cb0000000075ad177fa53827e2d0b2d93ab1e6b099c341864034009c13d5ae494352e6106d44bfde1e40f82fe0bc542154fd54365234bd13e0a0e4cbbf31, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h665d94550523110bbfd13d7f676262591a53baf25eb36351495c6f3c797d1d0b2a69f60f0d4a1277414a900c4eadc0b4, 384'hcd30032e93a773a2603955c040415bd3ba1ef4e43ab476dd4f6eee5825ed1bc5b0531099aea51909a51a8c6641e20c5b},
  '{235, 1'b1, 512'h6d22e20c000000000726c9469eebfd2e764c9b4750557869e51bef687b0b07862ad496e4c6a056d46f5d244f5f10ad0005ded39047ab8247ec969c4e42ec2219, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hdda8c851bc3920be100a4a1ff64f5415c969c2db653f3a8e62e950863aed9aa18a6cf9c98ed15725fba10d439ed94f3c, 384'h407f8f0121e96febb30502b28a64a8b86099d602f14ec25b68567481b7f42709c7cef8b212d23cd5c6fe7e5f00ecb2b9},
  '{236, 1'b1, 512'h5a5af3265a0000000025640fd363bfd88cc171f1966b1906138185d763f0ee7065ebd2a5813b79d02ca118763c60dcbda580f5ec322cdfb2c0a407e223f6b16d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h4c33b7661835f75c0b71e9a6084f58152e0067049e67732ea1bdf7788b1d5d7efe6768551a56f1633c6456caed18a5e8, 384'hf7b4bfcc041be40e5c24907c5174dd210e48725add92962fb223c1a0eaad11336c66612638a84b5865b50501f0667e9f},
  '{237, 1'b1, 512'h6c0f86f08b1e0000000069a0652407ab389f7f275bee385294bfc2a7a9119905f5ce4e1af41b3850d665c942f16914cf903717ff47c4e186c7fc97496a068b91, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2b1b1e7c87e0401be935919c509e020b391b4d5242df3584f465c316c88543a85f58dd7eca620e2c16d86068013892f5, 384'ha217fa8785fcbce6e5b1ad7d9bde09aa251a6e3e915df5f44ecb0d43baf33ec197537b2ac2d413663ff19c4d98943b07},
  '{238, 1'b1, 512'h5ab9d448ee67ff00000000baa93e38832a2709f7238f9bceb67b53fea917f665de9153c44b7280e1a5674dee745f5350bb3f2259ea084b398cff74d33bded951, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf3e8882f07c78c0b60915c078af978a79e9e9f64201ed51408e3776fd33830a06e6066dab7218df8cbafdbd7efeed866, 384'hea37a3525bd2b48991e3c82d8e9902693be65eb0953cb97a7f45381d4ba7598f9f076c0e4222c92a7d9dea7ba0668453},
  '{239, 1'b1, 512'ha1eaba175145939e000000007804c10bafa1416c6dc9d3311f844fe42868c6bdf283b946814df78822f198d26d886ed4713421a20dddcd82a21333d922eb39a2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8a37c7ba932e249987adc4b860a1447727b75d2396ae577e60a4333e116a88755b9b0bc9ab6f998042f455c5ca3efe45, 384'h2bab3f9a0fc3f0d84ad1fe4652160cb06a4776013741c5df39547534f53d255bae0fcec9a80b65b75b869616d798615f},
  '{240, 1'b1, 512'hb1fe8fe86f9994808c00000000f313a999ae7b5281bcacf933f05e4c8d526e761afa3141e9efefe959438620220c28bbad7047a6c1a98f95520baeb1d7af6278, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3dade5c9f3c3df658b91e73b5837161520c547fa930c0682e445c90a99ab81524200c3578703c815fc794c178ae113e7, 384'h866407b2dbc01d523df632447e01488ebf35a54944f4fb054cb89d31ed15bec3e8bceffe4a422ba27cb42675f37df5ac},
  '{241, 1'b1, 512'hfa3ef856182ec646db7300000000241a0e98fb88ce661de43bfd86f1c929391ee9ce6c05612b1609d6b8466a9c4d0af24ccb440f463cd18addf4674adb2f94ea, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0dbabe75fa6538e0861bbb502f930747fb57cb4dcd344db394714e0ccbba35ab832c42ad4895a0bae2148a4cd222f338, 384'hf46c223b0462a5dec8e180ed083736a86d05a29b5f1d600aef1b74bd37971d56d91661506c500260b5b51140336e66a9},
  '{242, 1'b1, 512'hed19e69c6f4de76b35ce6c00000000ad94175b8ad5f1fb69995d7d87abd893772b81ff83fd6caa25d1fe69b0317ec4068cdddac49512e6bf12d9cd8ce9a951c7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h810c6c1b6eed6396b6d23932a8dc5a73b7640c5f5af2af291fd867cd484a940ce4bf65f453c991e08d5e78c0eeabb08d, 384'h47920914c935727f8fbfe9ea3919998ba8455349199b34fc7dfd9a982bd686b08302171defc5bce02893c57a0d1b2737},
  '{243, 1'b1, 512'h2e2e984df4c5b45f7e337184000000000600f130d66940e8b4c0c1030e71fb8df7efce69100b9174baac3e7c474054e875f26cc182e925a17f55688964033e9b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb78c8f502aa5398aaf25ebafda69f36cf0420e40ef542d82e90e4a9a38ab4c7f35fb4ae418badebba8349e41aedf53c3, 384'he0df0dc985a24606c9be537ebaaf7dbda3ff7b0bcde19f0962cec1f43c42f2028187777693d08c07b1a9935cd1d1f512},
  '{244, 1'b1, 512'ha8f658c6632e4f474a6f1af1b9000000000048ac2a6121c8add714fb8cce854dbf1871b07a75008a42baa6cef01b4875eba4bc9327b41503cb36ac20f9354238, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'heebe681fb8e6ed44747d37513de1233130c99ee379610b6ed2dd389b223755e29e18184abf5a79195e202a61fdd938ac, 384'hc336c32e8342d3b4334369f49cc6d48e6d5913988cb3ac4d7debd07c4333a4612e2387f111d6c029aa65dc3cbfc5094a},
  '{245, 1'b1, 512'he89af705f005a4e1c5983824150000000094795c26507ca965c1eaf5782dd829a5fb5464eae46688a19ca7fe5851291f76fcd7f7226131d74cb4dde6063215e8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hedfaec6489e58021c699662c52fa0593bc278788380f3a5b13c42ff8f68b3e7afe266207589f331cf4a1e621b4fecef1, 384'h8fb91c6decd2d49c8d901a8ec43f7da91f87750abf72696d0c87c4258ae63ea3e5bdbc34e0031f95b36079d3791da027},
  '{246, 1'b1, 512'h9490ebaece67e31eca85b20871120000000077b2785e29958e0ab90faf8fcca953b142d51892ae5362246dc07a066ff6a4c9fed90a79fb59abdb7c8a888a9652, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hbd746ffa5059d9e887fab3be1c53c21d47e642cbd32bf3da4d1ef1e816e75cb02b14c58a6ecb50d4fce2bb86b8aa15fb, 384'hbfacd071541d1cec2cf97a82162aba7aac62120013a83514d7dcc35d11f5646bb1c00c3dc62b8ee74ac5688aa7d60523},
  '{247, 1'b1, 512'hdf22c290212fe9b66a9c65575e7be8000000002b9d4a3251cc7b64eeee3e76b7e65ac253a2e3d18658634eacb7494688a1616feaa0bf8a6cc0edbdeaa4533490, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hc42e5eeecfeb6f341a2c43e863bbc9bb9318e67c1464fbf0df53aee69156520a59c96fd4b2e833a531fd15e5b8a227b3, 384'hd9dad675a1edb4ee2f711177db77219d6e006572476a7d359baf2a846a3655a97fe2e4b109cf6b5dd4c7bc657df9a9a1},
  '{248, 1'b1, 512'hca6a7cd52432b20d8cc73c4e810dc325000000006ee638ed6bda85ccdf3b4606a300f2439910d382aa47f8e5839698e4bfa1756c5e93b3d6aee97edbc8ae7794, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf704c037bfc43538cea15d6fc20d034be90b0826ac65f64dfdff429c0ef0b84e96aaae207b2f9bb9eeab1d382d7634b4, 384'h7bed532df07a9f04fb7790836dd06e358388912d5cd7b5ebfdc7abd2e1510443297763d6a9460e3bb204f282a9e219d5},
  '{249, 1'b1, 512'hd912418a7d72e83ab66eed185bd627c70b00000000a88db442365b3ec21269abd09b4b2e040304518850835236add11fecca5a2c529f8bc4c06174a03b997830, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb36a254a2bec5f2dc62302457c20e8ee0747ec653b510bf9af9d9b9dc7ac05e4fd6578dfc6608019ad8034afd14da04b, 384'h73cdec3752fa0de71a3fa56e4dd89af0ecde8de54b39b638a1a3d85928a19e8c208feddf5d35a251d9b7350a4b183745},
  '{250, 1'b1, 512'hd8cdcf759b329e28b173d8582d7a91bb2d12000000001faab0678de44c1caaf5247d111c9e465596a89073d5492cadb0bc766620952c817f31a391f32fb27346, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h18dc650e8c186c04a7560467fe8d87eb61dff7ca400924dd3f36cab1c81f25281b69b18561bbdaab5715b997aa21c103, 384'ha65ab79877d06f7218f00ea72d871a77933ec8487a35f0ec21450567e6bd016d8878f36bc67655b4b09e8c765643e203},
  '{251, 1'b1, 512'h91f07f1a3d4b600628f1754ae5ec28d43554a40000000051e8c4594c5a2e68bf2f497bfbc7e703e1b18398a0b5515a38d60284b1a2dfad8c9132a7b9a98db6eb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he80439c807bdba93211dd1a63159b9a4dde1b627eec62f09939c0751cdeee9b58fa3aef507b96cd3ec819d7ac460c6d7, 384'hc0735ca53571c1601308dccf510a825eb6b959aed11cbfebce360c8f9f54e01f61b7195b07fdfdbeb5a4bf2b9af2d7b0},
  '{252, 1'b1, 512'hc6208a5a5c6b71a957477d8c39b01e072a65ac1b000000005c6ec3ddb8ce20911bba1864112d3407082c700820f8676037efb40be95619c9f686163a4d0cdc5e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hc673624116d7aa2943b60db72b9c59b734f937ea077788a581141539b0ddd3a82e4552cd9aed073cf234230dcc1a8e51, 384'ha4f93ed4b0afe9964565de3b73e77258a7ae5734564b74b8ccb1c7e612c2b4fc869237a6dfd317bbaf2bd75b08c4e678},
  '{253, 1'b1, 512'h7da7793b2bed3ce23ef7f1c04376791fa03f741f650000000008744fe10ac37fab4edf76492a339fe79e56ef75aee6c3169a0a61e3cb27e74666a4fe4184526c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2d9323897383e720a08d05f2ed51f4f4e267174893253fc6e475188f00ee881ef71fdfb19337f6800e492290b7b8a3e2, 384'hbdf5d45c4fb989db4353cca999065f9bfe51423bf61083b82b9c23bd2f25787f22ee5bcec9704fbb90a096e85dfd4cb5},
  '{254, 1'b1, 512'h48cd33f55583315ab2131d5db1f9cfcb0590b13a266700000000c9bd5d6fbcdf457e3bffd7b4875145a47be68b99a201b93b8685e80d61ce692a913be1183569, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7f31cbd14dbb0d079b43cca200e758acb429ab33eb8f99ad2c2e1f0be51d0e20e888bed0563f5d80a7ba603bc184bd52, 384'h572b79750ad421c43ca2eec7c73ba7ece9013c09dd02bf56db860ebb04b060a971d9ba043975abf340ba801ae0bfc722},
  '{255, 1'b1, 512'h1acaa001f6ed1b1a5b0bbde85513fe0b7aed266bd9da3100000000dc1113ab87ae3bf815157a1926b7bc3f659934702113570c26bf1bcdf1c8492f79614e844c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9c4559b076beb6a49a558d7d9bd68ad57f26c7d8f5b4a70a4b44182799810518e3ffa9e88e06e4e80792695cdf598dcb, 384'h977043d20870aca886b94b59d991f18167f9b846e64ce42c9c5f4e761a534fa178f99d8b9ff7d1d3119af4c206e3a9fb},
  '{256, 1'b1, 512'hc6244ad67598a847488d31d513fc9dbd21d96307c296a4170000000012f527d2192eacdb6045c48c250e317b7fc62ea79321783ae0f400ea4a60b48c2a2fc495, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h216fa858f98c2c36e1d63612d8e303ad1e79c2be9df56e4b914b39071e3cf6730519aec82e7a4b953387c5968c7ee2a6, 384'h9dbb30990b547dac6716a9663dec4adab95c8b9627eb82324960880c06652f95f2315f77963769be04baac725726ef4d},
  '{257, 1'b1, 512'h90f9b7739bb1699b90bfdf7cef079649e3f08242a08d05026100000000d3a4568eccd5ef4d94de4885986b68670617f552b9cb2a6eed337392b49ad4d04a9dad, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf4ade3885d93019dece7c2d0c60ed281e6df189389f6b32608d03e075f2c21038f6cdc1759b3121f4bcec62be0ced247, 384'hc523d6c83fdcc6fee5f250e801435c4bd6ff32702aa379f4e07634d29c5fc0c598a30332bd7ee235cf5e7cfaa121d63c},
  '{258, 1'b1, 512'ha7ee711aed6f375a8a15680f30deb6946501624b70b47c79d5a500000000ee6f7f0f2b69cde1a389e3abe86e51efe844c8e4ee7c3b2a15925d8c9b8b296ccc53, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3657272051a5892983150131cb07b1a10de3a82a366e2c18a630100e75281f77c074117a2bd0f86df722bdb779393520, 384'h656bf9b002f1de2a6a4e967d5bf2d1167594fb1e7f02fa8990d781568ee7986c2b161c3dfbd4e9c54b99af62d389e574},
  '{259, 1'b1, 512'h9583a32b620d5614a1c36e06ee45750fd69ef561faeecded2ff5b4000000007bb68b2b419fd574ffe1760fa0203fb1718c4e5d8a798563fdd98439f37a56dab7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0e6b00b7868ab7f1a7d738cf231f11a85e7df4c8b8e3fd0c64e3a261f986a20255bf60fa982cfd86fcbd6ab8769941d8, 384'h36b8107a327026b93ba8fc9d12c087ce06de3e7f02a513f520ba83481789a33a6667e4d96f54784b3cbe5f6133f76412},
  '{260, 1'b1, 512'hb6e404060dcf7182366941e77a0f0b43737232bbf9f73865863c271800000000a4ea51e31a92eede7497562eb5eff19b08310fdcd46cf3c22e069110aedc21a2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he999a6f89b37eb88add82ee5500fbfea4d085ea89aa87dc51a5e0231fb98e230e27cc7d8fb3f4cb50d731b2d9f95e4a7, 384'h684791d376261275ce5179bf38fd38adbfa0445855d25401566380f3ac47b97a5aa0134a06daeeef1b5cd1203b7fa020},
  '{261, 1'b1, 512'h57003aeb6ad8b84b54cdddb9243c65d8fd07ad1ffdd35f11c319f06394000000000aa9393490e8dcaf1c1e53ab5a7b2dfc0bd1dff4d0fc1e0c9dd5cbb035748e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h121df556b6e29fef7ccb875dc2bae65f8bd4b33621426d7fc7acc2003a016a95ae5fe3f22924019ef9e5f216bf21d606, 384'h97ea4126cb43ac8f1938ee82323c3e3177c09f8b7a7bb862fafc9cee1339e19329dc8a261cda1b050d782da06e79d68b},
  '{262, 1'b1, 512'hb47f61cf42394fa1c4c8cea80b83e366e30a938140f793851af87bd3782900000000d7a39fae605c98c96e0a5b0e8a58e47c3b50d4905171c884a64239fdd901, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hec2e792cfbc85f6e2519cfcd49e9b10e9f08a5cbe88a68c7affdd840ac21f053631912f62b3d45acb3cdf7db9f78f870, 384'h0a0da2d5e10886f7d4d7910ab6c4e589fa7e89ef94529320d3c6d168b8056af2b07b0afdfe2e3317618fe0aa1fbb213d},
  '{263, 1'b1, 512'hdfe80a6b887fa09cbdc8bb94300a4ad38f0380331a18c0a0b62708e590dd3800000000d364091041bb72f35391e792802f5c23fd676d0775e56ac2e41880d92d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0df1b7596ade29c09eb4a87290ec102f2bcba8731281a5b3818809510b2d3e23e0c2b194219be1144ae354512d4e4c14, 384'h710158c3e7816269bb08af3b8b1bbbbe595fd5ab77a06d14b47a9003f9bc5713e437135873e43c7014ef07ae8be2894c},
  '{264, 1'b1, 512'h16d0d407630fbd8dd9af18abdbdb902051c86b156254ecde6a5f0a5a1510f99400000000c202a44b1c172e1436f2252d80f9ab44794b22086f877c3bd4aa5fb3, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he364868bc629941f4aab4e8cb3bb876f396269d4f99e16eebcc5a8fe8ba787c2f226daa2990e1f6d5260bea7104fed06, 384'h99ad584fe5e7ad210592d5eb158a0cf28b19d2d9c74a688111367d254b71e39121f6bc1aa0d7f4861fe9f4d1cc2d9c31},
  '{265, 1'b1, 512'h519e4709f22b7ec44e321f4d403bdde7f532392786df003ecda243880f79f899f7000000000e3e6d749c0a602d959e0fd13a8a491554d233b9dcce6cac4ff3fa, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8e686e88746382c9371c8e779c271fcb05d10afa4b801bb45f9b48d35f2ef94a0859788104fc78b511c5324e209f658f, 384'hbeeec64ab193b195a2245391d51afd58a1139ec6edfee5a6c10a3ec9f71eee4caaf22d3df8931cca156fea6b3b79f67d},
  '{266, 1'b1, 512'h00ac9e66bf4db08b47a08e0b34e95e7ec2da8a82091479dabd2d57199b450dda70f8000000005b979f8077a5a74eaafe42ec70504f2bf8cd07aa23ef52c0321d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h11920756203720443ab0b6fd4f41788f7efe593ceb02ab61aa25caa1db7ba426e6c0719b44c44c581f14ae38bca2dc22, 384'hd6c6acaefab23ffe971cadad8386398bdd7bb986f225ef5c2f9c08cc7b74fbd679686ac02ca55c2a009f829fafe3c28e},
  '{267, 1'b1, 512'h2cd7eb20ee13fc351891dc4acccbc978161cc1b1e0cb95127485ff132176a972377cdb00000000add5eee3b407ef394da0255f21b9b8ca144d7e76fb075c6bc1, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h816f12f483675bdf87b82df29b287d2ce0bd281148c18ce3bd06b860447466164a8148d4db665d05a6fb733f7f7ba30f, 384'hda8e42ca2999d24b4ad0586fe9b85e0f78ca614a0acbc3c37a2ea75289f811aef84c9d6299737ea5e4cb1e743a2600bc},
  '{268, 1'b1, 512'hca402f2de7f990c5e1deee30d418810cd3a8707888fa5d54d3a5a0b3bab20144dbf37f52000000002a1f22f563f07cc9d066dfa8881777cdaf8a1ae4d43d6341, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1fd0fe36188f093ba2ecb8ddce12587583ea3638a07713a6f6573a9ffb4e50a3f6363fca961b8a0ac6a7f1414333f9e1, 384'h2ac94be5c224b12fb72375b22d52e3180b8a236b4980a6bae5aa4cb8119c54ab4cd89fc0682f564102517310e4eb2e1e},
  '{269, 1'b1, 512'h4386a89b56a955feed663fb88786a1c3916e8c65775648439638f2278c7d32c6d67f942e7d00000000d3a5ae2110db187684130f7aed62cb05159f8bb6eb1b26, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1e549378621758d1db17fd0cd84ec12031068c837afd13cc46cd8d0304230b45a544c7708b032505a048f627087e4703, 384'h261f1068011dfe1a99324e7d3fada3af75edddf3a84ff2d7089d587fdbf01a0a4cb49a6a1e8192cc16bb4cd37b909bb2},
  '{270, 1'b1, 512'h9a76ece71e15ffca113598c14654fea437156151bf5c8d47e15a6279ff965eedbe79fd4437f300000000148cc8ba720cd12a6cafa72448ec2cd6ad2852b2f703, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h90dcc3df567225a8ff08cd8f26921edbcab65e4996a6f324475ad04ce614c55adf31f568415be6f411e8b6ddb3252314, 384'h19542e3b7e26354ed7fea107c67932169fdd4f1d02d19ff7146306e93625ea81de67dac1686c7774a70a860feb8b08a4},
  '{271, 1'b1, 512'h24abce8b935764d6a61bf597db6c773145d5992485866070fe22cd0f6f871d53e72f6abbcac6ee00000000840dc44c1955185bfcf393a1786b04625904f03e85, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7cef758170e1aa6d553f1cb93f02e4578de16da89bb7434192ede200bf7c5f1b0c4c25e5e07ffe0889152d88cc951c79, 384'h673af79be286c8bc787a97af62dd06fc2e817489c2bcfaa9ef61b77a2e7b95c49af946cdc6fed8988ce4d502a7107187},
  '{272, 1'b1, 512'h3fa9e7c5fd635a7b587b56e19e8921e7cdc6d8f6b1ff03b579b907ccc2dba540c1782d5c35e3aeeb00000000a610ad03b540240313bbf54453b27d3794341d59, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h885c483933dc8b5609f0ebd2ed917b4820962db61101c8ec21e24851228f917e3e0bf3aed9eac628362b01fadcb88e33, 384'h4732acc7bf375d267f7f23fddc81c844fb23bc913b820ef00b23d0338a9b3142e20d93c25a22627ef78ecc22caa513ea},
  '{273, 1'b1, 512'h4025a46ad55fab109832d892d397d6e50c9c0aaf7136c275c259a6a61333a7e139b394a288148e32c200000000a3d26314f0694c5db5058ee34dfdd8fc2af9f2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7b990db18a20a82be2345511c7638c7f84cc75d679600d0de57861028eff93a4853d53c9d9779e7386ffc9f08c104d1d, 384'h17c38689a0dafbd6589558f87d73f1403d18ebc85e6ad071946a5aba27c9d833c12a825cf6331e5e698522a40c54c869},
  '{274, 1'b1, 512'h1e2fbff1179de8374cc3b5f47b00ade36b6494b8941aa810476c8b40e3ad3d7f5f60d8ff0d13bdc7683d000000005b2a7c0d9bb60d8af2267c656e800069cee8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h83f64e214381686f57693c04d640bf279a55446d3e8a43173263ab348b946a3b14dee892add49fa6057e91dc0391d7fa, 384'h84d489c507e32f88fbf8b8acd6fbfd3039da7e767a81d0b64a832f9d079c34275ee84a5cce67c0603df89bf36707e62b},
  '{275, 1'b1, 512'h1efc0d2c8682584f2504efc8fb5fd2848583ab11c97a1ad1d23db89d7d853316fd159eb4e2cee6ee4f2eae000000003ec9bbec801c26e55e61dbd6364bed8027, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6585681d741ed1019b408ce93408aeffeffb1888b3b5e0da5f2821bf15b168b2ec06a4a46edd8f9137c48480c08f13d5, 384'h87403a6bf1741ab398d49465ca99128740dae50cae3cbc66748268143a2f8fd5af0c6d727f320a81783696be6b642d1b},
  '{276, 1'b1, 512'he68fbb72e90ec509836476f39f26d3f65c5deffafd5b86448457438ee0c621fc8f97e83c77ecd131ff1e33e6000000007c2a942574c7da923726d5304e0de79f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hdf56c59e4b82d676c767e16c8c0adee66962ea6a8cd75f385cf44990257265b272e18fe19ca0573d829898bde3a33385, 384'h6ddcfaed53fedfc4d7ca7a6785dcd3992fa3ad6752c500ffeb18eb20c4a7994778f2dbe4ec1c827562e5100a5085fc44},
  '{277, 1'b1, 512'h90bc23f7e48f29ee5cf5bda8b42a6a8aed3cb6018636758be3051cee87758ed5998aad924516e34c49319b58cf00000000b7f0c29548e1c1244f0caff38b285b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h40fd073f877efa572a7e5186d02e1655e7e48be7f0461d7f71f218aa502a7d2dd61896379148efcf7ec30b3fb5943b7d, 384'h43cb9cf273cce2c30bcdc6f7825e4530687736340d01301050c858b4029aa5bbd24f08d56b07126ab48f74083e5d54e5},
  '{278, 1'b1, 512'h1c0e382d29f7ce824206c57f19794f9e8abe01e6af45a57dc9c01184c7b956aba27c6536c48c0951e2540bf566ac000000006db962ed4d45bf0d0c1c6c806b4c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h289f2782535cfbb90798dbc3a92434ec21c7f40022ab59fdb86f739dff5bca37b7a102db0a4f9209589e1dc88272458c, 384'h8337cfe11dc6b38ac8226b68bce4fb19f045f3b4c0da2185b49600176198509da073d9aaf1992e59640cb02fbd44530a},
  '{279, 1'b1, 512'h92cc3187d3326341d51f43165add210d496557c7a27669692c21c2912bc85d13d22a15ce9f2dc8052f89cdb3444fb400000000da250c8d1d81c198686e0c62d4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h487ee0974d8aed3ea9659822e128176faa5c576b4acbdcd2f21f23a6a13a8ee2829a88fb73ad332be5bfa6c2454a4fe1, 384'hea3b02f673a0c8f3144c1124b72ea9ffd2db4adda6210dca1408fe39028e3640a8395f73621315a47f505f7825e5de70},
  '{280, 1'b1, 512'h0ec91d81506646053327c352b11803f36a38ba32d940cdec35246744477eb4c423fd81dfe4e728bea623290a65646d9200000000f68a3961185e3a1eb3a74496, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h339911a1ac00fd099886425cf72263937cef82141558193a58f482b6e24abe1cfe5593771691da6b30246c7024c393f8, 384'h65a02c5ec22db3f9b8768dc7f5eefedc7c55ca68981eaf2ee0864477ac326d3e5038b97f059de1acb2ca3e0c369663e7},
  '{281, 1'b1, 512'h290ba1c9dd4ce7537613a8092317a721e35cf33f17d8c82bc20a765683871857d7a7f0f72e659928158b11760b339f16fa0000000065c91469026a04f6e368f6, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hda687f5087ea087b241f4d626f2d0230b7c02e66c0591ff642661856982c6939a47a502470deae8c69de091fe7eb9a68, 384'hc31d0283df38c098486ff90ca69787f1ff1ef59875db08d647bc454659fa84b9dac9834dedd81cd60bcefba2f945d4d0},
  '{282, 1'b1, 512'he9caa5454fd145db00275838ae34244a94ee61a025a174247c1b8056e6959c7f851f3038bc773457c88404c0dd497580644500000000719f683608f5718616e5, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'ha6bf038486ee5f960eb529e6e0e193a9bc2664017d577cf8167af1bc9ab079911aa965d8de11e352cbda6d7b4fc052d8, 384'h4d552856919ba4cf08ee1aeb0a3b2a56dc148a5030582a74317b39e1bb06e2539f2c978a5fc08fa0b9b362341532c393},
  '{283, 1'b1, 512'h1827524c50d2a178cca81cdd33a0be182f764450e04af569ce80811e55ddf11bf9b04675631ccc24d816b26e407df93f288bae0000000040fb10fffd72f8f6b7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h64d404bcc4d61394a7335d9a5fd9b360b07bea1f229045b803cff6847578dad242d1ccfe4765ba569013ed27da2f0715, 384'h05d970b9f318b56d86a2173b2ccd0aab2763b754098037943fb18ee1c5da8208cb545e81106d2354f563d8ef0da705b8},
  '{284, 1'b1, 512'ha5186acc06258c75ebd6c4985b00ae514a23405ece5e1c0a51122b5727c5b17a8adfca46c2479895b4121c304b5b2785c72c06a000000000ded1a008316d23dd, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he984af14b43e372cf258189a5c99d1b54e929eb929eb323da23496c6cc17a0ec7744ec97a712ce371285c23421528be3, 384'hcbdfe095d11e373cdf6b9e8b077bad25a549edd37c4e182f0b6b9ceb444c2e2b379dbce246466b6a0d764e3c4155cb4e},
  '{285, 1'b1, 512'haec77ef7d501e59ceb458f4b03194d730583d8282b6bb01ce0b0417143ca15c2059e8290afa26d6c1e38502d0b895bb4cb182dd4cb0000000097ca7caccc470f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7ddd669fc03d457c2c99b64a14799fcdc04e6ecbcb0c058f3d977e799a13677e6413e32737b39c3493977457236270be, 384'h386606a482a682efb740fd5df6c83903794a6708a793af7350623edd184ef61545991b5a06e121a66eeb934e972032f6},
  '{286, 1'b1, 512'hfac59bb2cb17756c53956cbb809fb1dcf8f30340a8b21f7a25a1e6b500284c29820250c5c8492ecb2f1c5906b55dfabfb8c47b418d50000000000efa79a0e20a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h68ac4b7ca89a38cae29905c9a535ea3311e3be2bab7ac1f65f95cc31627ceb428ef422874f1fb79ae42775d64c5533b6, 384'h6db4b6cfd5439fae0dc896332ec8fbcfddd5316bba8b0ea9b25a0bef8c3887f2f7bcd62ea2f75fc2ee6c8d4c1516842b},
  '{287, 1'b1, 512'he1942b44674c9c247d1f5857111e24baa87afe02ae74ac9d1ac122c10ced967b6243fd3055a4de1d50b98e24831c9f613d767a3060f7f600000000e5461279bb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h53cf0308ea4b28e52ce27123d6cfacf6e8deb01dde37b2e0f564b5587b30843cd8785f57cde322fdb9213faa07b5b484, 384'h8bcd5ad407f01b8cbdb18e42192feee4abcb231879cc183b8f5e6c888f57d48c2b5fab1d3c4369dbf0389febb6b3efa7},
  '{288, 1'b1, 512'h9ea149f211e7bd1f624b20fd50fd2c474d627b16250fb6281c6bf57af0b868f48101c656162b5e1415c87cbb7a685fd752937f97cf58a424000000009deec0f0, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he00f0b21a679d371878f3a4c924c68365426a98fe3e88c8d221be37ce5155b45a56108facf0c863066066f8898700c41, 384'h1fbe0b4096692ffa698565f3998b9bf8299d563ab54f4d0737e62a99d7cd4af970fa6918925d93b72518d5c6eb342c00},
  '{289, 1'b1, 512'he2d392cec1344167d947974fed90e637c5f80aba4fb00ba57dedea9f7ffd1b0404437d90e50f742cad5ed8b82bd136d13319934da1f04f50950000000059c93d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6697d087b2f535d80d744e3f36f1e6925dbfdcc91378a0da7c0a056e11458addc7cf822b3a2247589edb014615c9538f, 384'h718ebe1e4b46ace8e54209facf429bd1864e519af1cfedd58d9421eda697abc4e318152956a82876b1eaa41c186a72c2},
  '{290, 1'b1, 512'h40195fbc1bc4b600980e2c2b763857780d875bf68fa15558b038d9333a6c76f3aa4687e0325e29c3945bb8ac11ce675dff92bd5dcf0efe1264e900000000cdc7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'had49f1cda72a2d8b06a15252610a3582c999a9e7dcb0252a557c49edf42114d2fd81e6053d703415a256c2ab76862f78, 384'hba44945e707220de5cbdd4aff453ee42e8c98b17760fbc21bf7db7e85bb2461a69064bcf4667f00e3856d60208e83f6b},
  '{291, 1'b1, 512'hafc1cfa16e5549a03769a98e0a323b3ce3d8e3f316cd9f1007e4366b81a3affe3acb663d6a5d6a6857c736ce28eb85c432aad5ea98a80abb0b973c00000000b6, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h77f0603819b69683a871538d8654479e0f2e074a393ce153b9e192c94b21afd60bc093ec88373990880d422bf5d8270b, 384'hfb7e68ad7389276058da83963b5e544dccc4a61ad8b5377c42356ef6c853b363a3c4d8c5cbe93eb594a1ee2762dac2de},
  '{292, 1'b1, 512'he47ec71fc0cae21e08260f64fa9dc1a4c99ce92048144beeaf932a124c0f87a8b0db214e5424891f30a4cc0311efbb2d49807cc31733db9bd80f912800000000, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h77f635aba21e0010367e071ea7ba273fca770dfce16da8e2370f67c47e7096c33455e3a469dbe40d4ddb6aa98bfbdfe4, 384'h5109e7ebe6d89f80d5412bcddee586ffe658d08d18d34c3bf13af99e77d8b2ae265f32ae054d8e67053bdae80f1c8306},
  '{293, 1'b1, 512'hffffffff149aabbf287a78cde6477453f7f9c2310cd2d58ece43bb07019c69c965ca25e8df7696c97ee4ecd4966f7577eb41a60745d031a94f5856e1a5f95aa5, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hd9a417d59b5ce3079f364a9a04672989b7a22902d60cce65ee2ba15cd0ec8fd5191a16ec05574fb6119db4b639b9bc1e, 384'h85be5ab44b63d47cb215f2ccee2736af31e4d643a9ec43ba8d111f11758a6c7e73631031607de8e971a6c291c2fa6d46},
  '{294, 1'b1, 512'hd5ffffffffa5bd8691d54adc06abeae7d4857cd52aa3ebae84fb391361d804a381d15d6fabbedebceef14c94b5bbcf1560bc8b97cd4c4accead9b453f6d27746, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb2f6832448f8ed8107efd77c392d38f5997946d8bb47322d81276059bf0ad49632dbbee84ee0a5c3fd2598b4a262d906, 384'he2411b8ca995aa9711c2e273172c71d166fdd336bac39a3b3444c9dbfe9e3272486e4abf327eaf5b216bccc0900b7a15},
  '{295, 1'b1, 512'h9481ffffffff6e35dfab283e61e8f9a49de1cda44cdf1e2680292ded627b16d9b566ac057cef4c3380ee126c020a6ae86ded132faef613440c54185ed5986dcd, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hbce837f1423507353cdd93db53e9d468ff9f1a5ca680577441f222cf3c3b70931641a83b7eb18445bb55461ce842274e, 384'h797481a3380202e427659ba7113a5d02ed2bfdbdf88186c843aa8ed908956ee6e82eff7d7f1bb6dc2afb63665847d83f},
  '{296, 1'b1, 512'h2d8fbaffffffffb42e8498ddf2697ff4a2223fac0c486f05f57374d84dab9e8d13f52f6c898c8a7a74f2d48bee3cc16265e12a6dca3bee77c0ff0ee5e9af7e49, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'ha21859c29f1af1dd52dff9dee9ea6bba3e93411c2269a694e290fa6d47c10e6be33898c35880a9ebd89fd2795398592e, 384'h5fabca618898cfa105b61af5173a1cd9e0d9be0b15f82d2a31beff2b2df138720b80b3beef309ae980bd91511d45b446},
  '{297, 1'b1, 512'hae17b907ffffffff72c833830a0827c91ae711b1704754016d3b0ef4c8367a7e93d4ba6f63e6bb8d572c24bfdc55da0d39f5fc8def9b04723ae25c1b82a3ed86, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hc3490395cc64dfbaea1a75f147eafde602066e840722d1a5cf37765798e17afd531218c7db1d06e6fa5b7c00d11463c0, 384'h04626f800fc028ec0bc583c873bca0b47004f72d45705506b080747693e1f771966310d9c7031b6853047c936788f7eb},
  '{298, 1'b1, 512'ha55ecf9029ffffffff0b0266df6f2fc70941d6389583046c5649a1740aae64600c31269408a3fe8dc0975b57d60cc95053b7d311b677bda6e8a0d6792e328bb8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h2427377713b2ffcda16e539eb85d0f1d716ab5373bbc22c66d51789da2ff88c52824d45b260e0d1a151f0633ce62f483, 384'h0bee19617cbdf9001b57871cd486f9ddc0b022727d3508b59f9b465d6c43c17f101fead582fe99297f91eb9d4b552dab},
  '{299, 1'b1, 512'h37837a8407b6fffffffffac5686980dc2ad1a556be4d1fcf5dc000a18139c2322fb6d35995be1b96f942fa8bcb31b6d4c0efcdb2febaad183b00f4967c63c04c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf60077a94b71ab1d6a0547af84b53cc9b942a745644d14d16b17475030781cee1ba3976a55a2396c05b2e0c6afa13063, 384'h5fe9cf83ab2273b4115b5f55db9622b298424ed4ba84d6cdf89c1ee4e77d7799b874b47a53b51a5099b710939564ffae},
  '{300, 1'b1, 512'h148ae8a9d1f212ffffffff9007e49461386bac4123a9f847a6901d8d1508c822348ae29c100f38e169470e9a05b8cd6c780a06d49e062785dbdf1fd4cb89afbb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3dd186bd0227d623f977eb9cb66ee7542a555aa60c2d89d0d65b41def1201ced714890e3d8e9e5aec9a897d61b6803d7, 384'hccca9bc91b35e0a6eb86a3f89f0acd90fbad7cbdaaabc968a97cb3bde1f21e5e15809576afba10708024275a500fa903},
  '{301, 1'b1, 512'hc17991fc38743c0bffffffff12be8c0818873e8d65ea350547aa4cdc067cd0a4c21e1d9387ca3c60306f95160cc1f85a08ebdd4f3107b359483b719f5b9a18ab, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h5778c5f0cc38d1eaf74b185676ba2e7dbd1ddf2181402fec68795cdb66206aea6260289a77e1ab90ef29af55372ef2f1, 384'h95f2ed540f3e4c64b3c7f263faa36c557e5fbccfab96e8a0379486e642b579a0bc516aa8f58b22d0ca829c6b975d122d},
  '{302, 1'b1, 512'h45477dd24fb261b2dcffffffff376705fc972d1fc0eebc57960e96dbf0315340601ad9582193434f8cf1ff955cfa9a803a99d9465ab1d11337155273e65b2735, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h269baee7c333b24ebafc68a6b75cdc937be92337ab14985beed20222b7ab49b2db117d2622121202b42832450e6bb708, 384'hb030a6cfc43b6f2c431e93613c8104238bfa066a51d2a419b5ad852be40d69b63ccb2de9ab2ab0696d04f6a0058a8181},
  '{303, 1'b1, 512'he4d30dcc9e0b433fac32ffffffff83bb0169390c4443bfa7b7bc8a7c4421fb94a64d266b35ee622ee92a194a9c369a1bdd0961e4047a4fc3ed632b51f01547c1, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcbb128f0b17a20d422c3fa16f8889d1beb0f2e9c24b65719cc88a7a3ac51c94212daf1863814edcfbff14c05cb8b2998, 384'he826d9c348f9f52186e6ff5fe7dda8da26abc27a92734586a691a07f059558157d11afb316515d7dd9f1c23eefc13f29},
  '{304, 1'b1, 512'h8f46b06e493783b6d3209bffffffff5f263101ceb63bd0313945c63e59a123011230ea2a874c147574859882f49e6fdc842cbd97843daff440629f6a58573ee8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he51b03bf50a43ddb7a14524c336f2f8257d177b0a01557657a2e156a256ed8b0c75720b9e7fc5abaca512ffdf9a6d049, 384'hbecc64336b9aa348a9b3ed4ff09cf4f5dff27b730660031aec088858258d7caca3639e3d325311a139fca4c97138bc23},
  '{305, 1'b1, 512'h34de554e38945bbfefa7cde3ffffffff7b63c616e7853caa71db174d8c61626ec0c2d1fc20cbd176f51bd580fb3d6dbee8b1319ce824b44fd820e94589a562ad, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h177a00dce71c6811a3e303f42fbd84118106a28c65f270d534fbf6caf7af341b131c3dff2b9dab9732bfc13b8bcede15, 384'hb2b4fa6c519dcc3a1317e9b9f5635e9f8f352215c7066a8b2e5b953b1768c09f0e17981cce27d030b7f0826dfe468154},
  '{306, 1'b1, 512'hc80ad608a993f311fc5d85b14cffffffff76d81aa75f097430416ac8d6d4e8f80858d995030cfd10467787a708fb59252ba27fd5cb768e2b3cf03a351aec1402, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h9f180d741c934c8b5fef54986fe04e59c1121709ffccf9955eb529bb0d4f194cffae89079ec837aa71b36f6293b6577c, 384'h0e659e4149129c1ff578ef77fd645aa28bc76ef15e493dfda64e1c2130fa5936b45066e2678d7a6cb205c259140ceae2},
  '{307, 1'b1, 512'he9f4410a9857187394e0dbde1bc5ffffffff22ae4f317b16e8c82ca5e8ed1488b15705fcee61951d122b9603a8b3744eb429a850db99537b15bdee559ceb17b4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfd5d052c214815f462bf97f2648d9125d0b699f226879be26b581fe77bb060c2035daf878b2c41fbb1a2b59e91e91458, 384'h953d630e92a72dc4542389c31c07bb1acc4822a8d4d34989f1e412e288916adb8acddadaa903d0cf2528127b2071e26a},
  '{308, 1'b1, 512'hdbab4c37e253fc1deaa9e71c035737ffffffff6e927ee1da438de0d1d5152cd6d0549d2b8172bfeb94749da7ff020aa760407bc5e12a5a099a45a301588b62c4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hecd47c77cd0ad6d07b86e372ae85fcb26cbe86de5ea62e21265ec35df6912440c80252a0adb935de4657ce26d58baac0, 384'hcf1c88dfbe0782282ad26c38541e69376021ece2589f1fa7320c406bc8e32f6504e6a7801be5da4c5636887aa6dfaf81},
  '{309, 1'b1, 512'h2ad0f69e7f2e5efe8116b4b576a322e8ffffffffd986d354530161e2776001b50987f4eaccd1eaabb1c1d4d6c94e4f7460ebae1ff8cbf4a1df1cbf4a3e01348b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h415b96c16c2a4f837e429e5dd487dce404481e0922e214d4ca0952db08414f2747b6f75b8d8063f988961e34d343e920, 384'hda971ce9385c3dce1a36852482341f64f057803bbbb27e2f51f7ca6de19f818525a6206d9005ce09aea81625c5388394},
  '{310, 1'b1, 512'h69e08e9fa0546aec130be51f245d0daeddffffffffd8d24508cbc6106330bb7e4453fa88ddeeb7a8b80db338a7f66e078ffe0ee91d6b432c2d52b5a0a15f847a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8874629864ee14138b154be5bb497a0635554c7f21431222b29c169d702d27b3153e5503a32c68563098b8c336f5b314, 384'h46db1a0719623cd8bb38f15e3093ea829b9717f34a2219e03e0dedd9ae987d4389c370da97c709677787659f8996f613},
  '{311, 1'b1, 512'h21e7350eaa2b2a36fa211d7c6b144fc87b5cffffffff9c3a4d277dd4c34a428a3b35dc4d8c1840740df3876a387e6ae3c97b0a40325ae41007bb1de4338ded6d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb55460c9173b262db8e281a0106aa7ee28c41d6a3d1ab5eecad570ec32e9c41e8f98ff8f9818339f1233bca3e0f5cc2b, 384'h0ab47c58b0549a20e25e1e599f0d7c29a59869e630cb6e0ac559b8b7a330b197b396319439688131583f5d5992852f44},
  '{312, 1'b1, 512'hffde6b2d174d86702f3a46946c7167cabd18feffffffff2df58cb555aad0b0df043b0c01b91bf2ee4827aac1d987f3174e1fce7921c831a0b0aeab1ad1156fed, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h922662f604542fb01c35dbc904626c0c83883df72cc955589a82aae2305b50a57ca5c54b4ad3ce40bf49a297d343c22b, 384'hfb566679c426a12534fbe3fd28d60eba7b35a15256dba87e3874ad9851901963a381116394fce401ff87357fc18d4bdf},
  '{313, 1'b1, 512'h55260440dd65e8c48db54c801af143d639f08a95ffffffff9f03419e88a5145c37a3193cc07c160404a9b7d489aa324965d89fc40fab65a71fae34c56afa395b, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h7b1353d1112949c999386023a1f25fb63aa302c91846c94db05f462e372fdfab9fbef817fcb795e4ffea6928b1db9c31, 384'h0c1f69b6c15fef1e060ccf7d12f0ebf08202f4dc74ca1f2155f79bbf91bbff52984bfa2f396bb257d0d60f1963d7b542},
  '{314, 1'b1, 512'h16438d031fffee5b56365cb1a8f4bc19eb046a111dffffffffc16998d3235c27ddbfe7f1e45105d70ecb963cf511b0e09daa505bc426260466ec6528fd48b88f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h40eb566e887378be48ec5548a4974046fece281bf842c28067c781d10b1a64e83c8a1c0298d2abef720f523ab3b294a3, 384'h4f61d45339daa264848ef37f1d05f35b219df2fac7d0ac941790d4b7158b2cee19633d221193b05e1da473c39ff8d796},
  '{315, 1'b1, 512'hc0635b12b9164d0a9480ba133839afb60f79f6e7fa22fffffffff18d9363b5c503a5ae2f4cea06d8c5333965149a2cd0ed0491d1f9c8cfbf12fce9914dc22f30, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h88f12b559a6975c085118d3e2c587fc0706a2b5bd8faa325fac0e2ad3a305a1ae624ef3d0b59136e1ab6ab5137ea80b6, 384'h1049deeb0c9f6e6ce89efa749477b8c8b96e441c9ed0a650a8a2cd1f1ecfce9c9009b5ddffb1559d1a2dc40c71583139},
  '{316, 1'b1, 512'had86d31823a92384efee57d7fc747fc6347312c57d7e61ffffffffbad8263d3a80dcea096adc61333c39ceb1a06bc016fba8beaac8adc0692127ebdaf8bb65df, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h21cbc3b42183dbfbf11b1bf4852e358d8f3b3249c383d8f4d10915c37c70d8c77bca88f25ca18b2b30745d8b6e7b70f5, 384'h3e81a263ca654fcd926d9d21b4d0d95d0cb9c2a810d8d9b544c35805b8ae6aaffa71122ad28c0a6d4a7892e8392a5039},
  '{317, 1'b1, 512'h155ee257be62746434e431f20477a5a614b621ca050d7f78ffffffff517e6eeec93db0df6b6358b1f45efcb67e7b201fe4b0f7ef4fe49aed869621bb74d2604a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb651ad5599345c763cdab23fa4103e528b05602c8acf0121fc407000b3fa0dc6139f396472864bc203e1b5fc79281ba8, 384'hd7f573a9502e0f8bd7c6ce5511c21f16642fb81aa30fa4557f59cccf4a21b0c70b00b209413b28a0f4c8bed13b2f4c78},
  '{318, 1'b1, 512'hde8b1dea4af73e03d31712528653ece2fa048092693f2106acffffffffc4fbe785cc6cb125a5ca069dadd2dd809bc3c6246bc299c2bd84aaaef1085a561dd79a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h495ad55a38b11f61d891b4b771d180b81713c570877f5290b452d216aa6cfcddb5d2cbe63b14af2c83587aa128101538, 384'ha0c3586cc1585fc1a815b8b6d4b7468a0c3d493643768bd949af1e946439b9624c2a79a30731ad537d4c7a6638fa8245},
  '{319, 1'b1, 512'h372064a97724ffe3dec873aaa5c4e830fcd9ac84f1c4edb9a372ffffffff621efd798449ba3d7c009467fccb63c6e9a825df2926734122b80e8fc9a6c956351e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3560c7617e763a84e70e51790ee2ad764bab9f1f9701833cbe7daaad4776379140c71c9137b2df4df26834464b08992e, 384'hdae6f459e9df5cd64191a80e15a11b571d79ea08a0c0407355dd854b480ecdf22486881e2b3c632705828432817e4e56},
  '{320, 1'b1, 512'h0a55bcbb94c925c397b334ec37bd5216789d87fc6589738cdccee4ffffffffbca7bb2e94ddb13839ef8da502b39ac80f25abca143e0add021592ea7a36ce83ff, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hada0b173b36e55787f74d3d9e28c2464ea962f4320f70b568aa24119bf53056aa257006f1c375a5289c99293dbbc87d2, 384'h8e5bb37bb620539cf010082ca73bfb9c22244656eb2e1d846c2aac9ad2ef4473f7c702d1ee34d475d8c805a036b2d9ee},
  '{321, 1'b1, 512'hef503ce85b5b48ef35abff5d47345a71aa715f5e8e1568c9721a78ffffffffffe6124c567f2fb5b5f476271da455e079b655dc8c9506b65d9e3c60892984e8ba, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h918f44f0dfcbbe4f80abe5fd887f15f8cd9f6477ba38e5b6e367ab2b5999450bd06ca4653a9ddcde73804431db45002e, 384'hffb6be06f1f047e120aa347bb79eb41101881382dfdda5b7b25a87883faeb4f4f331e871ab075b259c1fd5c810bc4ea4},
  '{322, 1'b1, 512'h5f3afd4f98713d775d93b166838053fa503faf72cf3c00b3c57e0fe3ffffffff7b74af7667db987c9c205466e00679714af8467254f2e441ccbf1bdb9daad40a, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h4272a729473798dcbb582415bcac1d46b6b3b26510cab220408c964c9ed4499e85d3d45214830a256ad2c7644cd559a2, 384'h0c18795e6e2fefaf66e436c4ad48348752638cb7156eb51d081cc69cc1748a0ea555f924b1af8ddc89f2a07a25eb006f},
  '{323, 1'b1, 512'h9e670958749c5bbc0cacb1ee6c38e71eede821d75d84cc2fe1335af9f6ffffffff4e9613cec31f535c4c7bdab269d70a8d4b3bdffa3065d91435a4237cae96da, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he7fca6ecb733bc504e3ea6cf0f0d188233c4192bfd4738a254c12b3fe656b18e7e4432a58977decfd3e8a7a617fd48ca, 384'h4034834ef3566cb988cf77e544b49fc1194343bd1dbfc33a543b3e4eb13a004c4de8001d41d388ecdda6949dc72ad182},
  '{324, 1'b1, 512'h1e77a725c36046bc3bd6ca38747586093510952c0a3390d86b508479c0d6ffffffff25680ce9cd685ebae3cafde6315263f7cf4ea6117ccf870d42189ba3abb8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hf9124df58b5f0768b69a28ae0ba3fe953ce595ed662177795a7b82550002dcb9ad05459bd1c62832f68f464d5f67996b, 384'h68991ba84968923046726edf2386c7b0b09532e2ba04a424460106d2f3f55866be04d862eebfbfa186b61382452d8b44},
  '{325, 1'b1, 512'h59f9626626a34d5491d567d0315894fb702c1d7a2ec677a2b595a772b20d8effffffff20557e965f33f606242a59aea4cd565aecb931664e51fee93a92ccaab6, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h545c410f1ce821a1487a94f92226313693cbd1beee16f77c032449533b0b8d64cee954c31cfecc5f1b30b10f56c4becd, 384'h426b3126ced0b611fa37372f85fcfe3637479a151725c2d66500653a7acbd2c2f474c759e9434192c77c819135452b1f},
  '{326, 1'b1, 512'h001db8dc4aade36062b6ddb62bd342923f537cd35c957b47803909be234a3b58ffffffff0b537f24fbdbfbefce08b061b467fe60e7f86531ed3f54c6e29889dc, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8838a90a3b591c45780fb05f0546255ee9cac9a909be7bc3859378f11c0ce483db8a9e8cf3d18aa6fef99af08a47763f, 384'h53d55440575bd74805cb1af903e5ebe56aecdb51781f8386ecd5be528472dca4445ee4769faa6097ddc32857305ce32e},
  '{327, 1'b1, 512'ha05bf269c6959e1000f754963c2ee746346fac0d57bb119d3cecfa3dfe702fef2cffffffffddcffafb72da48023b4eae3593eb7c3c2d758c1c6c5e4dc57d53bc, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hec5bedca84cd99edafa98a82fe4464119e64d7c0ef8adbd314922cfb4f045e800e9e1b4c233d75eec58b0916966246c0, 384'hfe23ad017b4b525954b80b468566ba5f418e5e05782df4c0c8d2ca377bc7d9a076942eb2a3f2cf257bbb1e2a11642dad},
  '{328, 1'b1, 512'h9695a59c40d735b329f1f9c2ffd974ea8e66af6c65a1f7242e1eb02ea6721f9460ffffffffff9327209276e0633e07c96c9a2950a09411d1eabeda48ba90c8c3, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'ha686f038f8aba1e94cc210f2637adabb4f621a4da3015d424dd0cc06fd4049dff85b74fddfc6a84b7520c7796b7ae5fd, 384'hcdbfc125d7f03511c3316b5d3068a506c67645272610ff73b7874d8f4e9045f1bc9165ce9995f4e7d68f270659c52570},
  '{329, 1'b1, 512'h521abe64cfe7fa37251542760a99aba478c8b79a5eea4ba1fa859e6dd8bf23196e36ffffffff157c00247c6e0a683044034774f96f67cdea42afc9ebe8d78be0, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h88d55ac65133dab2ea64e7a30e35e8c8f8bd55636e4061e8e0dbef0b6052c671022c8c23c9225859ca2e72c7502f5e5f, 384'h8b08b7606d594f81e42456ad80062ba81d986e0ebbd3a0acb53629cd16112c84bc6b8e8949708271afd4407902684f5d},
  '{330, 1'b1, 512'h56f7dac71cfda3cdc27537a7fef1026211918d8041d79637eee4bf44f6fda371a67755ffffffff1dbdc9ce7d24880544364cd8cd5925c287a256383c78631a0c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1f478f2150092529b16a201fee978200c8c13c2b0f15e8e301a9c78d0ac8929b67cf8a8664e98e8caed1a0c5a856d8af, 384'hb1e546553d7efb04d03c7680e96fde773cb80207c8ec6b6d16db2d8b1ca3be228721694613d17801230e728bfea5370d},
  '{331, 1'b1, 512'hba44f1aa7dbd00300b9d114936943eb2585a2ca6cd8f11fd68794b5adabdcfec1919ade7ffffffff099e11a571237729c09fc81d86398317874c3722999b1875, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6474517a0b92fdc5d64e26e5d88616de83fc1be7e4ebb745575cd31cf04886fa07e00676b72e33ff6422e02a52b2d943, 384'h5a6c10b276d1fc9cd87797fd565f4a7b379835b16f4de07e4bcd4da5d5315943e74b5539683dc8e033249817b898aed9},
  '{332, 1'b1, 512'h125406f9b34e4f63c0a2288bf6166292074a0fed2b2c47822bb885520f2db3e2c58186b926ffffffffee3b259d2c85d9ab10b9f10f7f3cab27a8f528b4a82ad8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hbfbea37843a7008a368863f83d3b0994222d5a53cd7be1c0816e2b2e56fe50921e01729d938976250276b18f4afb18b5, 384'h940bbcdda97eb3e80715427a3b20df34ac1d293015c2cb46754a519ea6f81116f2c0ec780f81faf8bd3b35cf8564cf2b},
  '{333, 1'b1, 512'h46943ed052f77d2e9549dfb8b9a4c779959f7b0a78d6bf2dbde3be53634e232d52a793b7778affffffff162f29721e93b2c9de6629fffbe68596e94b26703923, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h925fbea8fe31438bc1c3208d848acc9416b2031e1a153fc9a25df2625d4a3e20c8ca045596d67ab3aff74add593e3897, 384'h878e3060a4b83f2d0a2e3d4317f35fb9fba0212e75e9913a26f02b35bd732255cb25d1db2910c1c18b0edc1696fb3c3a},
  '{334, 1'b1, 512'h2b88c2f7b3ffbf92cf6698268ef14cba56c268701a73b30436de1465b85a572363de2fbe10e2beffffffff9b6ad94f832c537e1e40dfd29f836574fecb7dd074, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h0624239416f6cf0755642ba9ae4aaf71842eaa1ed6e04c38c8e19909743b2660f0f191dbeecad3f2f53d8ef86e9c8603, 384'h87734389d9a063ca716f0915b5836c9ed840269dad20086eef59d278d7f13fd6748c0dc18ddd6953d6dcd9584be91178},
  '{335, 1'b1, 512'h4e29d13bd24e9f13d5e31ac769469a23d44278a67b110f7bab6095667a3a5180bc8124849e31af47ffffffff94e438c9abcb1301833210026c068417d2da4b20, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8037d7eb5c58311ce806a580fba2fbcd1db93466899ea527069812d41cfb29d0c092100efdbfb694ee6d5dfa1ffec274, 384'h459feded2c47bd44e021152160cd1e8be4efe37f6b96fbe79b9fb09d6a376023fa5f967a03bf9d3e82d3c30e9dc3cae1},
  '{336, 1'b1, 512'h5199a888f66bdde1285c6e1d75e11ca4a6fa67ceafbf32d81894eb60ba36c4786868dcb1384710d5d2ffffffff3d60d7798468aacd9f552c97fa4600343889c9, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h8f2dfef7d82610ab697f04ac6132dc2a5e5ac2b90db7620d7af3a58d8f66662c7d9178b39d87d187766f71a992c1003c, 384'he4e021d6d3951c25e786326191b47fb94d94b194f8c7ead99efe862d9f7d1256b8cf98ec671fc8b7b198aa91a16554e6},
  '{337, 1'b1, 512'h7692bad59be557b4e1db6cf148e5f0ff3c273d29d9017b90c8c26236cf78465b335a40716400ae0aaa34ffffffffd68ebefa85c403e0a25dbfeda3354bcc2a84, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6fa7a97e0a70f60703b691134e1d54708406f5f91c8dbc653ee953d139af4eccc83f565022eb109e20cb6aecec369751, 384'h54747ddb0d1ddab1b742596fa95468038e2ec102bcfa820fdbd324e4dc3c21e081259bf1248e591b38c5610b2fb3146c},
  '{338, 1'b1, 512'hadf9dc5a02f2bf38df234e566f0b5ae3c8b5a20cecc2f8565bb8f756ba59b295004e2ed1807a1e579596ffffffffffac7657366f92a09ca3685510feb2182e3e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hfbf953098613151d7dd1b4c949c71112f2579147d9abf50abf2a8bac0381f26d8bf5376a656b05a9d39c3a020dade6ca, 384'h1a3aa4c1547990302bd35a4bff0e5e85969f9ae4fb1faf0d7094149a0f4890f6420a6aa64a99906a6e4864a38077b764},
  '{339, 1'b1, 512'hf9db531c8bd06c7272a9ae2de6b4cac8e0281438eac5689c7f763241db7b88b4a6c71d53a3d03222f6195dffffffff0b690ef5a310f733b13a1bda4fe964a38e, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hc910fa2b3e62fa81ed99436a1954c6dca50019fe853e368ac4f2c836c8eaaa45d74cb2f3de1c492a5070cbb6fb00c94d, 384'hfee95b6e898dc053aa0426e2d0102c6841cb66ff0b43bc9acb71959d9e80ee4ab853a08900036ded7ebd9df3ca525e55},
  '{340, 1'b1, 512'h273f59b9ed631e0fc10467687508d817c2229d48e45efa2a6783290c6ab048c048a882eef2730e7456b3d4b6ffffffff0369568d9ede46d524123c6cdf78afb6, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h5c609212390b144969ce0cacd680d165422bb1dc28b98db296dc6eebe4e5dd84473e5cd901e416ba7f838b56b7af3611, 384'hcd1e77c240313a0ce8b4861ad2832fabf2585917d98aab7b2a525aa2f3394bd9214b930ce139555e04e51ffbba019dd8},
  '{341, 1'b1, 512'he6ded1492cb08b685e2c14f2f11d4bb2fe1601c47019cdd5bb3a42aadbb88f1335fe76ecf455cde30b30e18d35ffffffff921892b8870a2d1248dcd97ed5449f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb126bf96837a4bf7e09680f4c826e3ad4cb9edce04d2a547134a91523710ab99d45ad7de0c213c588a79db4a952ff5e1, 384'hc1c6ba25ea630772de4025689c178d78390aa50810c3ed17835d394bc4b1a568d1008abbfd1da87c0c4f7a284c77c052},
  '{342, 1'b1, 512'hef9ce8e0e84c667ba940ccb1d3317daddea8b9888a2ef5b718605aeff060c7140522f73cdb7670b0e055a2646509ffffffff81c895857965435d4c4421eaaee8, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1554c3cdb6a325689d85e7f1a97cafdc5d9d1586957c1be8e04b1cc3ac28a260f3c58dbaccabc3fdfef7cb344607be44, 384'h1259d8eb8b44ec7865d93edbdccc62d5f2d37e9f0bfe84219c2861d9bea7c7dd58e88c2f2fc14cc586269a28070010a8},
  '{343, 1'b1, 512'h388b354799942c6595ba49bc6bf8e7ca5c06c6ae8015c0f58e69192d96cc60e30696c1284ba98c1b22c5c7f23bf8e0ffffffff15f579e355c7258262f0fdfdfb, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hed2dd0845ab8621992c4507468586173d00ccca7faed06913db70eca582667437c6f589be97e5ea5c6a0065d593a3cee, 384'h9016b1626e66fe53b5a7dd6661660b2fd735995b1d64d914c5c5c6a91452e050617314b14d57e464381c2730b879414b},
  '{344, 1'b1, 512'hc6bf307fea8c2799ef482911ac86779072e5757f934a3671ad8c5a9e372bb2ec8d318ee3bd0cc4460f9050c937a3409cffffffff81c81c22e9468fd07ec09f55, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h58a36f6b0ad5a0211d5f58e2f74c7e7930cdb7efbbf45d0111ef606c253b4bd227a7e53c834619503d11113582ccf013, 384'hcedecc59dd9f3ece325fde05c09f0e20614c79fce3996c71b5ab2b26451e832b476b8dff9c8a67b655d8499a171f5e71},
  '{345, 1'b1, 512'hf5f21b002be6b7b3a605b3bcc5a3a12aa0b905565d958028fb8c44d8e5182b6ea4beafe63cbdd96daef63b98ae46ff91bfffffffff3ffcdb29cde67329851fd7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h217e55870cdeb394b937e0ebca9cceff3d1d69ef2c0f4ccec8cf95b912d544caa244b1233d5e677de94c6a59048562d9, 384'hb716db65e62fcc5f01426ef316ba17c612e0e5d3539e06a962211831f118cb0beb10f289f32d7ff276f119c234359822},
  '{346, 1'b1, 512'hd88d68932ee321d611334d87de84ef4240025f9d0c8f11bd9aaea2e7729ad87ab0ee66d229b2eb78221050b375a54bd698a2ffffffff0967dbcb983a8f09417c, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hb2bc708b7e0616f4b1128cd39397554cd046218a7385198f9f52c62ba10431eba1cc81409ae6695f7e29d7a19716aa87, 384'h1f34499351f6d29d222e08dc498985cc7230d4e7f49c2070b787ae2083e328a808ffcb047d89bc0e2bb295a6f8419f4d},
  '{347, 1'b1, 512'h611df311628ef69305da2acf952b7289eaabbf389dae756f08c459819db39b7133f02dd126e0442f19bce8ee83cbaabdcd974cffffffffb7195ff14e2d445864, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'he2d36ace4a4a5aba6c06afcb98fde61ab464d36c5f52fb51b9678e76bfc6e8bb131b8a118fe5ddab580a9300d84602e8, 384'h1ce43e58f9f03d52df5720e3cacc7a46eaeacda51d0701581637da10233a0bf28fbacfb411dacbda9172cbe4b1b093c5},
  '{348, 1'b1, 512'h4f34828f9520f17da9e588884a26df5ab85e8456184bb19001abc926a180c32a112ba4164e81d69b8fdaaf3c60619a7d1a5840b6ffffffff8748db5ab09c4a64, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h3f3357cc7dfe35a0268195bfd14187fde860a12f776978a12a2ca43dc0237bc48f475bd440fdcd43ec101f4d552bfdd6, 384'h68555a3e46b373adf3464329d392fbda0cb3f2490c7e6482c888755f62aca75ed416cd59bc0f84fcbc749af79e145d64},
  '{349, 1'b1, 512'h4a3d25b54b17b001046f323462e30475caa0fe686e8fa4eaa3b0cbf604de9812e2cb4eafbbe44222356c1e1702c09078e7df08dc98ffffffffff06067e01ce41, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h26bdc539d084e97356bbca9aa23b52ebfe99fe6d26027b4252cfccbc9359cdaa4a526faf9ffcdc0f831e338baf9bdaea, 384'hbce39066652e0e83c85affbbb56234788f1466770d9d81f014e7aad4694c167f06ee3bd0644f983415256bea8274540e},
  '{350, 1'b1, 512'h6a763ddd1f348cae57162f918abd67d536a03431ed29721e179403366c3fe64f1083d4a64cb7a9fddc7c5a3487675be4078be3b484ffffffff2d5a70dd12c49f, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'ha977c3fef54b995745c8d34b56429b8deb9ed266a2a782b80f954afdcad3642bd1ac554c17d45ea5d35038524c960f8d, 384'h21e318cde939f7cbb2fc842b0885acb3af4905bd07a834678f8229e74f3d3d6b779f7253cbf0b1295da1775a43e956f4},
  '{351, 1'b1, 512'h0844602883dbcf60972c8b943b5ea020ccb0d19c82eb86cb18d4225a79f97279539214d6e3df6ba6af165c9cd95b8b67a36b39bbd101ffffffff5a9aa9794dd2, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h80f7b25aea62a1f244dd0b4938e3be40a5077c278e0624561b9dc71c6e530557a8e362ebb5e7ea5244b06d68d9862118, 384'h5a7f8b1dce45583bd9b9dd6b441126bc21526ce861181d2eed7a4bf9998ad4c6461da3107b0ed05711f744236f4d5d9f},
  '{352, 1'b1, 512'h73672c1037e14e2ed10a0928e8938944667e83879d16f2688f2fe0087494b9f496471dd4e27f5cfddfc4b5efc4e7fcd511d2f67ea879f2ffffffffaebc4501e4, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcb33c16745d056d2f5450f88f77f10f27a405b4e2fa94d9dd71efefedae568723c036026d8911d987bf43f96ad726a1b, 384'hc00433bcf5a4d87f937fb8b3235ef87e525352164de2f28f96d332022e8437b0b56c7eb3a28cda7f71c6661fe8368ddc},
  '{353, 1'b1, 512'h1c28cbb7dcfe2b79763ccf8ebcb7939ea373f7751d8b3965fdcd8b62e8360f619321855d0fe872fcbb3509f48c195d96b1d765983c695686ffffffff51d7cbd7, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hcf6cf760e836a2bbd6d355890a6c2c342196a39d2b6e57fbb8d01ded5639fe5d2c0291074d44758cceafb816c3a1687d, 384'ha1ff948964717d567b54d8c866f79ec0e6d147f7e5dbd6e266efc3c71cf6b6c116a6c2d675f1664520e8775545f7a056},
  '{354, 1'b1, 512'h823e30e3f8bce86e5790d073d931eed5a7ab1f52fdaa4a2522831c73dff05fdcc91829a51c8c0c97c24def713b52643ab17a700ddfa0988740ffffffffca2992, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'hff679d0731ed5aa6973a29dc14e56ec983521c0070600034acb6b845b9c01bb3e01bd86974495f70a919bc8991b96023, 384'hd68741cf8770abc4dddf74089cab8679cdc77a807f587f6b112dd8fb7df47c469d440bedad5f3615e667c0e0689e66f8},
  '{355, 1'b1, 512'hf2104bf641a8b485448e73c4b7de7fc4ec1d3e06eae0f264dbdadb0d514a7aa2ff1567a80e8156c2bd97579eb1467c0efacf0fdd1166e87838a2ffffffffc8e9, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h1f42b6c6ef17ec124bfeabdbc78fbc18b3773d7f3001719bf83547aed7bd8b85596d39c3d74ed5e39e558f2367b8c5fb, 384'h0e42b5d0addf488e15881d80abcd4710cd1cef8138fd41e868f6edbaf369807246b43e3d98e141a7fb34f25c8d8f52c3},
  '{356, 1'b1, 512'h3db47a2cad8a1c43f31ee677cef231cda0f3853901676c1732771602ccdcc294a38fb8df77d5e6e5737d4c8e05953aeb81edb39a25931717b3c154ffffffff9d, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h6aecc2ac6bb44f69f328f2d26ceaaa8b92fbbffcaef5258b9915311afc47259ac6cc03e1a88211a603c7342f0fe24706, 384'hcdacb0fcb3c54d33420fd48331c5db26e4bfca9b7465c9b16163d9ec75175442d8a37564ea372d57a47a5828d8ccbcb3},
  '{357, 1'b1, 512'h6becb022ae22ffc4efd852cec1259abcbd9936403db48920bab66dff9bd34bd1ba5c30d1e8752af80d13d9304dfb864e834181cff7e8be9467cc3617ffffffff, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h834a374b3ec9b7859bb08427e9d880875af3c1a98ead009f24bab9ebe1d067a13f83fb78705ee8ac32e6950fc7a2aba4, 384'h43949adf582e52ceefe9e3ed95a0c4a228da95705da24102b93c45b09fa08ff9d358d98f8cb681f68434485695c43909},
  '{358, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h2da57dda1089276a543f9ffdac0bff0d976cad71eb7280e7d9bfd9fee4bdb2f20f47ff888274389772d98cc5752138aa, 384'h4b6d054d69dcf3e25ec49df870715e34883b1836197d76f8ad962e78f6571bbc7407b0d6091f9e4d88f014274406174f, 384'h87658b9215c91a52e1b82d92d9ffd6cfebefe6433b5c46cfbde751da58b2d44b22c2da1dcbbdc9d0d606c53cde2d2ffb, 384'h89d6a04210e58032c0768adcd13120835cb0fae97d1f387e4009df9154e9365f1788ffdcf854bf7b9eea893b7f397f01},
  '{359, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h0b478a0cbf5eb4671e50812f1945e4f852d8890dacb40e9947ab238e6db8f1f97f0ef769e44a1c9455ca0f21f8cc24be, 384'h4b4b3e825064d3ea8bf8562e7a23c9a61026f77251acb12478d3391e5b08f9ed5979b2ecb974d5025b683f146f30dc3c, 384'h000000000000000000000000000000000000000000000000389cb27e0bc8d21fa7e5f24cb74f58851313e696333ad68b, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52970},
  '{360, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h0b478a0cbf5eb4671e50812f1945e4f852d8890dacb40e9947ab238e6db8f1f97f0ef769e44a1c9455ca0f21f8cc24be, 384'h4b4b3e825064d3ea8bf8562e7a23c9a61026f77251acb12478d3391e5b08f9ed5979b2ecb974d5025b683f146f30dc3c, 384'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffeffffffff0000000000000000fffffffe, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52970},
  '{361, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h8482baecb7ce217056f34fc8a85875876002bba5e13fbe9857d3653aa30f6821d687f5eb4a2be7ff2c0b29a2e053abd9, 384'h0d3f5d116ce9307f9f6016d46ea72bb29eb4778a0480b1dff8f5ddaf458c788c16d3ee41398b72cc7b5c60d811517cae, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52972, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52971},
  '{362, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hd71539a7304a82f93aa69f89f0668fa273dfeebd1ead07171de49f3d071d5dc53a130c14d2189b8c032cc915a83422e8, 384'h8023068f0154419b434a9ce0bf12c99235595f4b616c2db97b28e523f947451198fa63aa7901e71f8d9b31bfd2cf7ad0, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hd1aee55fdc2a716ba2fabcb57020b72e539bf05c7902f98e105bf83d4cc10c2a159a3cf7e01d749d2205f4da6bd8fcf1},
  '{363, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h0f2ae91fdc85f7739a400be4c128dcfb377559c936bdeee620cd08449b7bcbef992c2534dc559cfe328067fc3e87df8c, 384'heca1b61fd631c99bdeedc28c4a780d10ab38fca2cc7ed53eab34309646d5c2c9dc7063fe5a7a58426e66b0ca3db1c22f, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hb6b681dc484f4f020fd3f7e626d88edc6ded1b382ef3e143d60887b51394260832d4d8f2ef70458f9fa90e38c2e19e4f},
  '{364, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h1718de897c6b650a9c9212a0c0e67a4698e63c3567f025e6e02dda9161ece01ea0a18afc29487a5ed01a48856c9aab4b, 384'h5e4bacf9f45d4659438dc28ca21a0c461e38cbf911471e4141630f0f7c32d4aa7a1310d48eea3a413bf682201fed3f27, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{365, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h93f92e69558939a64304de24eaf2799ffb29e3dfe00a8aa354317138c2942d449fa735eb5b5ec24429b03194fde99240, 384'h19437f8818df2d550f0079f98571c83b75ac0ca26edd24793d0a95068d8258e17830763b03334ffc8bf5476488a7c1b0, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002},
  '{366, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h969e39e9e2f3e48996e7faca4cc842790f8a1477d1c5699933563b470495f4ac68b76d7e1d4c39a7b70df2dfec1a0816, 384'hf03e95c8b98c478330ae3e15e1b80e33caa3057f4305e84865d3a270cab9751214947d0bee6a23d412d19e606a9839d3, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003},
  '{367, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h969e39e9e2f3e48996e7faca4cc842790f8a1477d1c5699933563b470495f4ac68b76d7e1d4c39a7b70df2dfec1a0816, 384'hf03e95c8b98c478330ae3e15e1b80e33caa3057f4305e84865d3a270cab9751214947d0bee6a23d412d19e606a9839d3, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc52975, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003},
  '{368, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hf9feeef209b372bb678d2d1275c653d7bdb6908982879321e7f4ec7a083ad85762ee1b9d85c7227bdfbc56e44727030f, 384'h4c57fa58b619384165a3b50a62c63dd3a8caedc6204cd35c404d1f16a6cbbe8283228448b468fdbb12d54e5d2cd70cea, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accd7fffa},
  '{369, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h20d23d3e5a68e72896db6b2500f0797de558586f31d79b696b19a170299674024dc8acb4adbfa2ea83b0e5deda5adc8a, 384'h20534957096a651f2ad6ecda4188496639d04ded5039df67b3e7d28586082007021284e8e11f79bedb42cb5a7267e55a, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100, 384'h489122448912244891224489122448912244891224489122347ce79bc437f4d071aaa92c7d6c882ae8734dc18cb0d553},
  '{370, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h5f662a2de99ba5d6ba9d441581b1e0036056dc2d8a146080fe4cdbefa47efbcda2874ecfa49f4f8fa99ac309d917bf28, 384'h3a4117e5bc5014c832fa8e08eedca6c642d6181475151c1808b3e33fcfd0103a1e4210fbe8ff58355f8f6706743e0cda, 384'h00000000000000000000000000000000000000000000000000000000000000000000000000000000002d9b4d347952cd, 384'hce751512561b6f57c75342848a3ff98ccf9c3f0219b6b68d00449e6c971a85d2e2ce73554b59219d54d2083b46327351},
  '{371, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h22c42feccc69d4aacb408ba1d1f114bf54c90489792d2814b264248dbed9e156a64835c9ea97b837120d2a717f584841, 384'h2a50bb39dfef060efd1a6dfb23018e7601d3b3ba80f19aab9e334cd5e1a7db144ef25d3745ef40099a510fdfb837070a, 384'h00000000000000000000000000000000000000000000000000000000000000000000001033e67e37b32b445580bf4efb, 384'h2ad52ad52ad52ad52ad52ad52ad52ad52ad52ad52ad52ad5215c51b320e460542f9cc38968ccdf4263684004eb79a452},
  '{372, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h9dac20d645bb55d57cab932da900871184be9f92057aabef5af11fa2dc0a795566ee35d94b00ddb3a0c9d09e522a2440, 384'h9681ec7ec2a90696e49aabff89fd7bff27d7a779b3169000046f0566bc14580feb9e3a13b0b045970e13e58265a0be87, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100, 384'h77a172dfe37a2c53f0b92ab60f0a8f085f49dbfd930719d6f9e587ea68ae57cb49cd35a88cf8c6acec02f057a3807a5b},
  '{373, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h715a3ddb84b71d5921e96b1323d2d129e7c1fa16e31c0ebcea6b233ac8cfb61258875a364f1d3a548f09facbd001709d, 384'h8e03bc73a762cf14f5470c8fee9f9650e7f9d808b1c81264eb9f85c6e94bff9ea398a88a0b173da4b585e0eed4352cb0, 384'h0000000000000000000000000000000000000000000000000000000000000000000000062522bbd3ecbe7c39e93e7c24, 384'h77a172dfe37a2c53f0b92ab60f0a8f085f49dbfd930719d6f9e587ea68ae57cb49cd35a88cf8c6acec02f057a3807a5b},
  '{374, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h36d3a9ed200de6c6ebb1efee2d3c30e5f72c521c57a387979d1aa772d57088764033bd9da81bb73f8e834eb305b9444c, 384'hc8a0b783cd1999ba35091372ce47e096b6e29ea54386f7501d7a7ceca2978fa0b3b3be95e03f883c27b38bdc251af860, 384'hffffffffffffffffffffffffffffffffffffffffffffffffc7634d81f4372ddf581a0db248b0a77aecec196accc528f3, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{375, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h31a7e388c243a6dcc6509df7ba5ecc2566db33ba6f71d494140daf8fe0ba490859cf9d524d83eb76a06c02d616f508ab, 384'h27a272ac157f661e1c0e9ba5944943d3e102bed4c52ffca7232cd8b955e0e792d982a7fa849d9c06ca1442354e1b3171, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001},
  '{376, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h31a7e388c243a6dcc6509df7ba5ecc2566db33ba6f71d494140daf8fe0ba490859cf9d524d83eb76a06c02d616f508ab, 384'h27a272ac157f661e1c0e9ba5944943d3e102bed4c52ffca7232cd8b955e0e792d982a7fa849d9c06ca1442354e1b3171, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // s=0
  '{377, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h7381fbdb53668ef60581152058fe6fc0fd38605253fb9b9d58e240893e8da5ba4488e5af092f431b5a359c4ac62a67d7, 384'he75d552ec90e3b6921ae1347f7609ebfe1524eae34671f824261ba3455908102be99e0231f929c718fa970286156760b, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{378, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h5b896e18f0747794790cd9155c74d60bf5e9cf6b34b5c43b0776de78745c2a49414b24fb036e5ec658d00f0b5ee7af8e, 384'haa7569743b2c97130e6a92cf9c74c090275f09c4b7299f3e38c6a559bdf7b75cd78b291b714b4f2ae1b25878bc005608, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9},
  '{379, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h0db3126187c353c0034e618ba3f4630e0b706312ec5211b1ac91f01caa23bee17456b5914e10c5cc5b9decbe078fd3c7, 384'ha332aa70d7486cc7924ed61ec8a1b045ceba0f0a55a4bd3e7a9497dfbb1afc7193b6a34a8c0f6bf4dc5c707df14732eb, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294b9, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294ba},
  '{380, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h0d0c15cb6cd38bea588f92c654f2c5b36d3fe1db8cae4f69dcdbeb51084e0ccadeb17990c1be62a55a32ff8df78157d0, 384'h90ba4770b1f1f2105fe3ed29fb793aaf6fe220c630b4fefa096460eccb31153f1dc6696f650d95e85681f229f30727f7, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed28},
  '{381, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'he3d48751eb34c96700557036cc7cbf49dba0b6761c5f82dfe122951aed52045612ec97f4a1fdef3105bf720051bf0c78, 384'h8fb468400d982bd9dbdf9a44b1f383eafc6420da722788085a5745baa750164628c1d7e7b7525fbbdd93d9308ef49ae9, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'hcbd2518ae59c5c357e7630cbd4c4cb1555da9a1d381d9ede05a3783e9fef3c1bb2aa85d6b0a80a5a6062306811743c4b},
  '{382, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h8f326a3e9ee7e1d0927439d925cefeb8e1165029930ba125c309788adfd1dec07834392ec8f8cbcbd8f217e203082d0d, 384'h5b6d713a80d496832e65d75936d4407524470b5f74304b075ea9484d18537af60054e620bd44fe4570a7bfe4242e9252, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{383, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h289ad7ccd69eac6bb4f5f104fa8832159c25fdbedc2dc0e010bfb408923f5e22cd7c78886e1d1918a7fcdb04bcc1dcc5, 384'ha0e14f606516353edcd0ec7a0be00da3bbeb465fae7af639ee01472977b898db57543460a46b3f9044f812194622b59e, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'haaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa84ecde56a2cf73ea3abc092185cb1a51f34810f1ddd8c64d},
  '{384, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h93fdc301fd5497c6bdf34008e44b544a4491c53fd03e68f730f2e0a8a696665425a6e18efaa72add19d7040f6daea9fc, 384'h021ebf043a0dbe24c71741975a45f15991aa0376bfeef5c7dec3c5121f98a464097ede93dab4e46205a4932677d52d86, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h66b9e4d1b3768bee2b2defbc0e6911a38e0c774b97f62060830bb641c2d50a8ba9d8872f4ae86c33d327562482b20789},
  '{385, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h60cca8bb9e1bfaa97a3be18893c7043a77712deee44b913c939ee4b9601157feb515208125fc7655e0fb359307e0cc3f, 384'ha4e53d3e06bd1002a2678182a95189c4890fe6ff1d4ed9759f4690ca373a766fbe4caaf69f85d696ac6745da022fc5f7, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hd3aacc47d028c849c7635156b94bc4aeab9eb29ccaf794fc0261569f9c8912ef6266ed43956849a2e4c0badaf2edc39b},
  '{386, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hf5f7dafb7cb762f4a86d038828add9f5a1bcb59421aaffe01f5b2b7009acc3a097ac12b792b149c36878f8e0fd9ff441, 384'hdb91e4fee136dbd5d7f2404a42d9548c2edfeefde40af2262fa1e52553485c9ff689f3820d8f075387225e782077d485, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hf265d814894ace80d5706d12daf316f3450758b9c581286b807c89fd36449c04baef8ebe2bc988825696a1470589a52e},
  '{387, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h84481d7dba583052bcd1586c4a99f3e21b4eb9df66381981c8343289d28052a2d50b41932d209b93c7ac3540b595b048, 384'h1b6b0510ae966673280f1f7d12d5a66a2c69762c50821c191e93e906fa4ec44588ae8fe8f1769660308268f5df019f1f, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hcbeff5c13e09b437cbd2518ae59c5c357e7630cbd4c4cb1528c147efee6b14dcbc0fafcf1c116dfa4ddd7a042a79da3b},
  '{388, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hbe352e662168556652a4e25acbb593c3898d323ed4c9dfb00fbeed0fd57601d910d226facf06c13b64203f21a6c1f8d0, 384'hcbbdb29fd0413bd92f9376ee5848b90be84fa9b1d5eb5e699120036fd5c6df0d721e39752fb01848a3721c01c3631981, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hff5c13e09b437cbd2518ae59c5c357e7630cbd4c4cb1555d71296100da3347dc5f026c06dbe99486ef3463ca655d88a6},
  '{389, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'he1eb96d55fc336b196fee593d9d42e0c52ed45ab2a90d9a07724f6efbd4d51263d2f6e1d8450ede4aee61a86bb7c0ae8, 384'h8c5b22c8c7bd73177963dcac910f2f184131b7968914bddcae43812bd3b66a7aeeedcfccacf02b9854b81c1d54ef98da, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hfeb827c13686f97a4a315cb38b86afcec6197a989962aabb1aef747fc02f61d965eaca5b6f228192f17cae29fdf5e7d9},
  '{390, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hb5a2e0ded857a339984938bb7eb311939814a1671bb161bd45fe14e441ff29535e84b6e6a1355176b2d4c90cfa063a57, 384'hdebcd15e16b32a5aa86597310da1b106d8882d9967ff4d58f1dfb4d77c58aec4582ca97f845a2bdcbb200c6f6cbb09c5, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h3e09b437cbd2518ae59c5c357e7630cbd4c4cb1555da9a1d2a658646e12f71ed983b89459ac429062d11f6ce0b53b14d},
  '{391, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h29e5a700b55ed124ce61db14feb891c75df37797b96d7430b42c0dbc0347acd6dfee873d9eabce23a64ab3bdf7293103, 384'h254b4fe4502daeb1d261f33ecf1a87e81c19d1fcb3d6c4147e2fbd2fad21ef25a8cbc641809f3505f9a148f65adf694d, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hea4d0322e1725250d3a21591af916a45be6105ed6e774b0857fbaba69943dc1f411d9b1c1fb66d2b4b722c09dd32e210},
  '{392, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hf88f95de4285d8e1222bb900aebefc42d7639a9c4af0baed4462e050d5395773d8605d3eb7ee3d9ad9c29bf9a50e33e0, 384'h43b63c509f022c7752d18b255834ed0b282d2a06b7587f7838fec43346d686b255742f460eef623d48ce2da5129f53f1, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hfac83b5ab08fa2d2263f04e12ee07ab55562a902ec02f649340351c805632f4bc78ee682b97c97c47877e884207044ef},
  '{393, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h58e9de6249a28ee74438064f2c57a5b04139d13d1fe310399c64e886d7817798d88aa6e8017724457fd67b1444271a39, 384'hb7233c886c537589a6ec877a6140a85926168b2bed502c568810833d47e5a55b6410be70feab39791fb4277f347adbc1, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h99461b2e4c897411d4d21043f196ee5c71f388b46809df9f4457974031622353ae418682fdc83b4719c4c3464a1321ea},
  '{394, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'ha6734ac30bdba9498dea41492041fbfe95b3359c2cad630d4e31d1c0a10cba666738f35de5b7ceb56fd29c08cb5611da, 384'haed6a6876ca0e33b7887ea0964681ef703e861337493ebf6d54ce8db740ad207c755668f89dacc36edeae1a5c0036a05, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'he5e928c572ce2e1abf3b1865ea62658aaaed4d0e9c0ecf6ee68362e04a1334fd856249c47cac58eaa6a724e96f1cb2df},
  '{395, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h45db79275eefb11d4a0febe14b31c1fb6cc4c6a0aaefabe674ac673e09cc844499d8fda96ce46c59fa43ecb8d3cd115e, 384'h9116df7b21f6e27e53e6fb2abcb37586f22bdcf02cd5c235d71e083240538079d39ad7946b48d808e32235536a89f58a, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h7932ec0a44a567406ab836896d798b79a283ac5ce2c09435c03e44fe9b224e025d77c75f15e4c4412b4b50a382c4d297},
  '{396, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h185b65203c076b524d888a491a6e934a33b1fa51e6b7ee5fa3a304f9c1f08991ffb3d4485ebdf0f984b0f45a6ba7e149, 384'h1599239305c4d9f4cef234ecc6000bfd3d771969a7671d4304b0ec1a1a6154bbe26d99a57b1c5e75e1b5eef7447a8fce, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffed2119d5fc12649fc808af3b6d9037d3a44eb32399970dd0},
  '{397, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h58502135c1ced850e12947e2702f4048dede7754d6bef88cb599eb65fb326af1a4008540d682c21ec1469c9fe4801e42, 384'h88df3893083bdc8824ba709d4247f8a29d1b5135bc11bb42445f4f6d22821024a7cc7975f475a0d5022682855d7c0ab8, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h79b95c013b0472de04d8faeec3b779c39fe729ea84fb554cd091c7178c2f054eabbc62c3e1cfbac2c2e69d7aa45d9072},
  '{398, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'heae29d829ad084552675196c6f394556fbd73c7e10a48b8620282d4d3896ee0ab4d09996916c4ddc53a7cd3c3606d3e0, 384'hba37a1bc6db922bdd12c34c5d9478016d4d6793ede0aa18bb491564460d2db30c4016e36839ba636fdb908bc54468156, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hbfd40d0caa4d9d42381f3d72a25683f52b03a1ed96fb72d03f08dcb9a8bc8f23c1a459deab03bcd39396c0d1e9053c81},
  '{399, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hbc31a5f5793a1a3d81bf6dd37a55b13624081691990a5737645ebbe5a8f3921c9eaac0f23b9174c88451eb61c69d0cb8, 384'h83bba1948e818dbba902f5e184a534854c69c881b85f682ac12dc019e1c6d2da742bfccbefc5ed84e95b42930c09fc50, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h4c7d219db9af94ce7fffffffffffffffffffffffffffffffef15cf1058c8d8ba1e634c4122db95ec1facd4bb13ebf09a},
  '{400, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hc76cbc996421f5acc36e665635759cdd2d615b4a497bea9c321fded0cbcd3546c8ecb7ab587b9fa4fd5bde6add66ef68, 384'h7ecafe0f227b59c452ee3c77670ad9bfb8b0373821d8c08821ccfcdc6f1938efa612e98411f99f50279f794b59e2b10e, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hd219db9af94ce7ffffffffffffffffffffffffffffffffffd189bdb6d9ef7be8504ca374756ea5b8f15e44067d209b9b},
  '{401, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hef73af0706ca2030f3b64d23172f6f961fdad25e7b68151b81e59fcb0b46a297786360b85042e69bdb4c21c189d3ff35, 384'h892c292dcbd50e19905a9b558ee7f441ad00130c7578e13b07831fa13859610c7408974e3b2f42e33c9db2436df40e89, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'ha433b735f299cfffffffffffffffffffffffffffffffffffdbb02debbfa7c9f1487f3936a22ca3f6f5d06ea22d7c0dc3},
  '{402, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hecbe4a557d3ae0adaff67f90c5c3b46541fc570954e00487af5e13c9df150807feb76a38ce9a4dd11f847f8db79ed97e, 384'hdeade0c36705e4f117d02ea0966e0fa01d0a31168899cebd32e544dae19bd59486cb10bac77ad90739c1b3a8744076f0, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hb9af94ce7fffffffffffffffffffffffffffffffffffffffd6efeefc876c9f23217b443c80637ef939e911219f96c179},
  '{403, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h3be024650ba1e28f3b6ffbbbb7b2fd932d97d966b576c9fa2829147787225d3bebcf6fdf52ceceaa97f3e713321ae05b, 384'h5202ae4f52a80ae69dbba2a647f0cdee63f132ca4d2a56180e1304b6ea49b800e368380696fca50d2555bb8467010a9a, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'ha276276276276276276276276276276276276276276276273d7228d4f84b769be0fd57b97e4c1ebcae9a5f635e80e9df},
  '{404, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hdf85a11bb0c9c5f6a4e18b3ddffc6c597fd68319494847fe0034ff8aa1b9df00935d617ebb69d2e6524a856df4333b62, 384'h231fa6392ec16aa1ec13d144777c6ad0264cbb5020744d1bcf43f4d1c3ad6962d0d41c1f62dc0ba1f36f3d8b5e72e670, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h73333333333333333333333333333333333333333333333316e4d9f42d4eca22df403a0c578b86f0a9a93fe89995c7ed},
  '{405, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h6efba105b9e276b04ecf896e141ff172027b1bbb18bab6c29c1db29dcfe7a912fbb28feac2346371811b79a03459e19d, 384'hb04f05153092410e09f8b52da437051112e951d982862e0a5ea61e8c41a407db2d00a7289d3531193ab37f6f8ef4e7b5, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h7fffffffffffffffffffffffffffffffffffffffffffffffda4233abf824c93f90115e76db206fa7489d6647332e1ba3},
  '{406, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'ha82be5ec5f9deed5ca6d104480abb903ca317671e76e232a900ee2bf2474b097ade520837168a4ed5cec6dbfcc0ea0ff, 384'hbbf3498d2b5fe438b2ff9f450c0f6db2c20c63ca120278f97cc8c188afa653914a6e40fc9299c578e1d27453eaf77e0c, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'h3fffffffffffffffffffffffffffffffffffffffffffffffe3b1a6c0fa1b96efac0d06d9245853bd76760cb5666294bb},
  '{407, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h45a99ab80d9721656e0097ec2929fb96318e99759e1559fc754e74c6d240ff1495ac899ef6f6c1f434e39eff0cbabfa0, 384'h05c6b0f31de5b9bfa20ea28a9070a6f3322908d5b0bfc0d7d3a8cdfa9e93b653b4768b454011beff9bb9bbb838162bc9, 384'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 384'hdfea06865526cea11c0f9eb9512b41fa9581d0f6cb7db9680336151dce79de818cdf33c879da322740416d1e5ae532fa},
  '{408, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hbd44171238bd66df3d410669d961fdcd4cf0d635f30ca6a3e4228053ef0aacaa24cb55890945ec5a57f3e8ff21cfb542, 384'h766fa8a382f21dff2c3803018c94b52ecd28b7ee04f76297026ab13707ff68afd98b39d431c46b13ef3cea81b4158770, 384'hb37699e0d518a4d370dbdaaaea3788850fa03f8186d1f78fdfbae6540aa670b31c8ada0fff3e737bd69520560fe0ce60, 384'h213963af02bb080baaa19382bc09cc2ec5d8692eaecd7a5b0fe49250ea46ebe897ff62811de1980ee73b0e4354a15e62},
  '{409, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hbd44171238bd66df3d410669d961fdcd4cf0d635f30ca6a3e4228053ef0aacaa24cb55890945ec5a57f3e8ff21cfb542, 384'h8990575c7d0de200d3c7fcfe736b4ad132d74811fb089d68fd954ec8f800974f2674c62ace3b94ec10c3157f4bea788f, 384'hb37699e0d518a4d370dbdaaaea3788850fa03f8186d1f78fdfbae6540aa670b31c8ada0fff3e737bd69520560fe0ce60, 384'h213963af02bb080baaa19382bc09cc2ec5d8692eaecd7a5b0fe49250ea46ebe897ff62811de1980ee73b0e4354a15e62},
  '{410, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'he3be38a2438036a73738ebc1babd703a9d001b681f069ba101037e5874cbf49b9aa5a0e114e89ad7135bc0975d47c891, 384'hc206de0358a77eda6b6c8ebd0ba5af1d3fe8ff1d8e18841a9ed9adaa7c13d430531e36311a559a680f0fe7afaa7fa2fe, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{411, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h33a24f4337d8a02e4a1ac37befe6ec55169baecd409cb75e2980281d07cc12081de5d8602be39dddd1a2281785b15c32, 384'h9e9dc79417c0ea1958b9ec8073ce60eb159f6aec9762496ff0416013d14d77de9c9bd215b396253704195aaa2e5ad174, 384'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 384'h33333333333333333333333333333333333333333333333327e0a919fda4a2c644d202bd41bcee4bc8fc05155c276eb0},  // OUT_OF_RANGE r_len=49 s_len=48
  '{412, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hbcc18cbc9dadb319cbb464a6bf13c3fc23ffe396295e0c6629d6d423a95a55e9962d95bac76e5cec92be75f7400becd7, 384'h01d4032a396acd89fd62df36ca522bbf580a870f65d40eac8b734a1e645873f554888ae17e69c61bb0e0c85d38fbb78f, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326, 384'h33333333333333333333333333333333333333333333333327e0a919fda4a2c644d202bd41bcee4bc8fc05155c276eb0},
  '{413, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h3674230033c5da4bba115c351cf4544b97c76800938af5d76d1393ee2541b5d318c305d6f3f60fbd4840cd3e357b43b6, 384'h9f79b78bce247f5800af3504797cc14b15d5d4213106b5c7ab83e4a7d5f6dff31ecc12ab18caaad8c02ebb234215bd30, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{414, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hac7d897288e85320e94487ec773f2e9c421657227e742dfc9068273826bcad1a9aef4bc63ea74d112ecab091e5139209, 384'h7e797b58408de6b5f9adb46ec302e9e373887934e5a79ff5db51188b997cd250935b505662b66abcc726be81446bccea, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{415, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h6ccf7c5d5a5ca8223535dcb03823673058c686cd9560ed2c094f3ede52dd0de59e5edfcfb829b0a95f939234c931c361, 384'hb06d1b75f60f6c9de67548dcf100b77e6a667d7b6bec104a1cb86bfd4398127ce9ed50a3756ef7cbafb68c01e37349f1, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h6666666666666666666666666666666666666666666666664fc15233fb49458c89a4057a8379dc9791f80a2ab84edd61},
  '{416, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h5aea5b66a22e9ad05ed948050b7478d66d52bf5c8ae1b037bd35dbe36f90651068b929e294bad3852877f9ed8b56084c, 384'h88c0ff92b7bbe5a36cad9a31baf4a8da756e7b13169d1b2c2177e0c119c91ceddd8414a5d29d862f12bf1816636514d4, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h99999999999999999999999999999999999999999999999977a1fb4df8ede852ce760837c536cae35af40f4014764c12},
  '{417, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h4dfca708a087c8165edcc21010dbc83890e895a61bca93ebb32913b7c1bab5f13794978c0a8f437f9a193f3d49e87c99, 384'h968d673558b512e86a3c04557cda68deff647165226ecde4a53eff3b3036e88259982cda28365608064d14e7d067740b, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'hdb6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6aae76701acc1950894a89e068772d8b281eef136f8a8fef5},
  '{418, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h07dc1276082eabff63a3b967d64157e68d8ae79491ae90d43a79c1548ce1cbfb48088e2b256ee8a4d6466d676eb82a3d, 384'h14566877ffa534182760363c94cab0d4ad8d3a3fac2d78b98dc65f8a78b5484696a534d0894a029e70cdcbc1c6ce2e54, 384'h08d999057ba3d2d969260045c55b97f089025959a6f434d651d207d19fb96e9e4fe0e86ebe0e64f85b96a9c75295df61, 384'h0eb10e5ab95f2f26a40700b1300fb8c3e754d5c453d9384ecce1daa38135a48a0a96c24efc2a76d00bde1d7aeedf7f6a},
  '{419, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'ha82306a028e2fb16f5b6eaf6fc96d3430104486a35d25a35e66522a5f68f53e4c6def3893009acd8c75abbdcdd93acf5, 384'hb6eada815252a46fd996d0fe4a735493cdea3a0a9f617ff9469df8c1b64ce2d95fd132ef398de3014263e95fed4fb213, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h55555555555555555555555555555555555555555555555542766f2b5167b9f51d5e0490c2e58d28f9a40878eeec6326},
  '{420, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hb425811b3bc72bac8bb8b031e9d9c36c550a70dad6e5245e22f0b8c42c56f0a628419d04f3e89879f261ccf1006af569, 384'hec26b6d4eee78d11140e5bf311e7dc4def75f1cbde623bc2a5462d50cb478b61e9dcca74777cf260bc8ef8b7cdad5e08, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{421, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h5b031a8020ddb66a43f05f3085e333101f5fbac8737a867f6e83efd108cb2caeefd1210494bdf774c788eec1be43d606, 384'h19a6290c3ccef1dcb3bac46556460254f5079f43bd5470d366770bdd9048c3c3109b67438adcb965d6a695d2a16335d2, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h6666666666666666666666666666666666666666666666664fc15233fb49458c89a4057a8379dc9791f80a2ab84edd61},
  '{422, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'he17bc4a1caa870988f63da22635337513f59c055fb7dc873eba0df125dff66485d87bef520ebd4c576c0adf37db80d5b, 384'ha6f702b447a50c9fc3cc87dd0f6d9a1707b5ebcb80dd3c0bf891bdedb1f235ab33c3f3e4ef7334e384a24efd503a0924, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h99999999999999999999999999999999999999999999999977a1fb4df8ede852ce760837c536cae35af40f4014764c12},
  '{423, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h051590a4cbe93ae21dc6f272d5376b240e229117b35f9cb892fb6a7ee00c567eb5b7e951af15251733fbf83e3b4a2ca0, 384'haf4e5197d271ad16eb6561c186013a577bd17f399bfa20c908237c7a784d5fc3dd98665f20f85fecaf53ac79ec7f0017, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'hdb6db6db6db6db6db6db6db6db6db6db6db6db6db6db6db6aae76701acc1950894a89e068772d8b281eef136f8a8fef5},
  '{424, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'hc1d95813b50699453f6b4859f2ea93c6e48dd46ea154786afa5f01a9ea7093761114885711285ed7bf78a66ad0f5fcec, 384'h09342a946ef35fd9eada444687903f43640025cd2a1c2ca4dac580ed933d9fa9441ad80f3ae76b531acd8abbd4d672aa, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h0eb10e5ab95f2f26a40700b1300fb8c3e754d5c453d9384ecce1daa38135a48a0a96c24efc2a76d00bde1d7aeedf7f6a},
  '{425, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h3617de4a96262c6f5d9e98bf9292dc29f8f41dbd289a147ce9da3113b5f0b8c00a60b1ce1d7e819d7a431d7c90ea0e5f, 384'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed28, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{426, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'h3617de4a96262c6f5d9e98bf9292dc29f8f41dbd289a147ce9da3113b5f0b8c00a60b1ce1d7e819d7a431d7c90ea0e5f, 384'hcbd2518ae59c5c357e7630cbd4c4cb1555da9a1d381d9ede05a3783e9fef3c1bb2aa85d6b0a80a5a6062306811743c4b, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{427, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'hc9e821b569d9d390a26167406d6d23d6070be242d765eb831625ceec4a0f473ef59f4e30e2817e6285bce2846f15f1a0, 384'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed28, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{428, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'haa87ca22be8b05378eb1c71ef320ad746e1d3b628ba79b9859f741e082542a385502f25dbf55296c3a545e3872760ab7, 384'hc9e821b569d9d390a26167406d6d23d6070be242d765eb831625ceec4a0f473ef59f4e30e2817e6285bce2846f15f1a0, 384'hcbd2518ae59c5c357e7630cbd4c4cb1555da9a1d381d9ede05a3783e9fef3c1bb2aa85d6b0a80a5a6062306811743c4b, 384'h2492492492492492492492492492492492492492492492491c7be680477598d6c3716fabc13dcec86afd2833d41c2a7e},
  '{429, 1'b1, 512'ha69f73cca23a9ac5c8b567dc185a756e97c982164fe25859e0d1dcc1475c80a615b2123af1f5f94c11e3e9402c3ac558f500199d95b6d3e301758586281dcd26, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h9404b3ea09d8e0777f2f492c3f15736ff0e63e22389c676f9a1463b8d8153bbce5e522ee992cbd8d5e3f9378d33969fa, 384'h41593e5eb1eef51f034ee2e6384d17f5f466089bf064567571839bab3ec4cfb1a1b8533011e7cc3f9e337865385f86f1},
  '{430, 1'b1, 512'h86fe1b4ea7ac8e339d04e40087534c61e245dd4a0c22754a0622642bba56de900b2d431e859a36b1a5ff71aee560522eb0d3251e018c2cb6a10b82031cfd37f2, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h5662c815b9d1680cb027cbede73cbe0281b02fa97f99e6070ebc442d90dace4a8e2dc0f365c149bda35ca473e920cfcc, 384'h367cf31980d9dbc7ff6a0a72c1fedf525a29fa3e83021f387030bc465607d5e65aa31385be28c2000b6a01dd83c8c02b},
  '{431, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h4a886d736f5b9cad6044bc73f6a753af24c68ec366459f4d6bf9bddec936c8ee913e4c88490dee78ebb7234ea44b221d, 384'h67e53c5c9a53ac2879502e4cc6bb16e896ca89b931f439aaf91e3bd9686bc01d171eae952975ed2e8e9ccc9492fea51f},
  '{432, 1'b1, 512'h7d795fe6a97761d89b35f64e09555951f6ec2a669a9fa03481c100ae158f183e2171e142437d2c3a42352108a22a7e3d797beaf6c3075db419b6f4acca479c83, 384'h29bdb76d5fa741bfd70233cb3a66cc7d44beb3b0663d92a8136650478bcefb61ef182e155a54345a5e8e5e88f064e5bc, 384'h9a525ab7f764dad3dae1468c2b419f3b62b9ba917d5e8c4fb1ec47404a3fc76474b2713081be9db4c00e043ada9fc4a3, 384'h458766812c6e6818d9c26659700ff3d5f9de570275d0bb8faf16e2e28990486288d09b825424e67a738a4917dfb1afdd, 384'h9383ea7a3b618018c1dd12c5df505ea4191638746578dcd700c086c6bc132ea028090eed26a7d4b0ffa779081fe3befc},
  '{433, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 384'hacbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'ha4d7ca043122dc46bda79650f5e1872e27cd9aa89744dc897af249521db2292650fd1cd66cebff3a3650414b5e1a70e1, 384'h7ad031bc876682105cdaeba7405df3684aecf89586b63578acd005b5b61360c9e8cba3a8287a39fc6322138f962fda1e},
  '{434, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 384'hacbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'h9a8e7c526acb3d0be87cf359fa1c7fde02baf47dfbdb4b48a2b6814346f3dcdbb9530a652873739d9493b807046f8d62, 384'h1c5781b742217b9465ce9daaabf6f94d4763bf362654092f9f23a8114b840229201e978353ce9f70a03a78f537967a37},
  '{435, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hffffffffaa63f1a239ac70197c6ebfcea5756dc012123f82c51fa874d66028be00e976a1080606737cc75c40bdfe4aac, 384'hacbd85389088a62a6398384c22b52d492f23f46e4a27a4724ad55551da5c483438095a247cb0c3378f1f52c3425ff9f1, 384'h6bbb20407a282269df53e14e38f4ec8075726a93dd2623f3b947592e57cb26f1d306ed79f02512d2b926ab0d1e8912ff, 384'h6789df1a3e41a6abbddc319e864aa536df09a0d49651b65b7b1a4374dec51cee619103ed202b22da0e223034299f0ccd},
  '{436, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hd1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 384'hc6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h5b87f6174fe9312c2c9100ebdee5b3c8ef5c33c03b2a2056eaad4eed7e0634e73e62b2ff5653e880d1bf2a5ecb165a95, 384'hba21de53b2c2c925688088358a4997f4a2d9abc98a46dbf1277fc3221107519c2f7acbd13ddb13bc9bf9130e680378b0},
  '{437, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hd1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 384'hc6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h2fba05c6a994859807662dbbb5b7d09b1cf70bdf05578636fc8a19d3f887c572a26027fa21e9f7831867f414ecdd27f4, 384'h73cca8521906f6aad663b7def79e8ac0065f1c74c2be117b43302981abd47083226f297c7ba5c7b93ef359670cacff34},
  '{438, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hd1827fc6f6f12f21992c5a409a0653b121d2ef02b2b0ab01a9161ce956280740b1e356b255701b0a6ddc9ec2ca8a9422, 384'hc6ed5d2ced8d8ab7560fa5bb88c738e74541883d8a2b1c0e2ba7e36d030fc4d9bfb8b22f24db897ebac49dd400000000, 384'h41119aedab871dc7a6d2dd8bcf56e7d5297d61fd422096d550812a0d495a20d7f6765b733cf2e6c7c74a38051c71ffbb, 384'h11b37e5c0fbeecbb4ae1f390f80c3dadea079e7a1bc0ca3eb7b5b09fe9d74e1aa0557b0ddce29f0a15f67781ad2a671b},
  '{439, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 384'he6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 384'h2cccd76c899e528e85d6a310b93ea35113d3feb569246818f3b56bd3b75dc7246fa95cd051416593a09094c62a946e48, 384'h6d305b01bd4be2c7f855ee71c2da5cbf97dbb8fc23f6a887b8a365aaf1913213947ed4a07e1ead5741516e13eb70b64c},
  '{440, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 384'he6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 384'hfdb90442feea49f2800a28d90f18421068b806ca6d088bec08bfa3df4fb7e866101d92e294d6e8b98f2efb52e57c8fe5, 384'h351f5065b69f2aa540d50e551965fb8a05bfabe9a4670682aef61a5ace5d5fd9310ab4a5b05f9c02f375ce0b5b6bd8ca},
  '{441, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'h1099bb45100f55f5a85cca3de2b3bd5e250f4f6fad6631a3156c2e52a33d7d615dd279f79f8b4baff7c713ac00000000, 384'he6c9b736a8929f2ed7be0c753a54cbb48b8469e0411eaf93a4a82459ba0b681bba8f5fb383b4906d4901a3303e2f1557, 384'hc183e7b548dcf2668e7414cf5fbb82c0158d3ac4e76a7862807682d954a0816482a601e6b6ddf728899bc6187774bc09, 384'h529f8b1e60c9f641f380a3f0aa39ed7eef7828a943c977a2562a41eeff040b871d422b9b5661d12d605f963eb0574f6f},
  '{442, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'h000000002b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 384'hd1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'h7a29d180b75d661776ed0e5d0a720792a88b5429e8d6961465d5bcc871094141441c37b996cd0f9fd05a1b42210648fe, 384'he4a559272307a37bca803ba8306bdd42bc8fd1e62e21df178c7f9ac35003d05ccf303885a48c3fc8c8d2bc1677c8f00a},
  '{443, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'h000000002b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 384'hd1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'had44bafd37a9f20b1c273fc604f61ec68759d956c47d25787d74925b54ad8d32f95ad49d1f6eaa847cc1fbb405008df7, 384'h3b903e998f4d28156dd66e7954fb10d2a5a7f1f70e8402177cddf5577737bf633909b3037080acc469fb6ae5f0b33ec4},
  '{444, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'h000000002b089edd754169010145f263f334fc167cc19dae8225970ae19cc8cb7ec73593d6a465c370f5478b0e539d69, 384'hd1951d597b56a67345acb25809581f07cd0eb78d9538a3f8a65f300e68a1eb78507df76de650e8f8ee63a5f0c5687c98, 384'h7a2fa750719b0b3a342a7256fb4e274a3783da3569fcd6442e3452f35bd57cb669fc9f93500839a2b76c37a986ef6cb8, 384'h34d8ea62222b7c3b71b776c322d2be021621fad3aca0a1cccfbb1f390ed171158a0919e5454cad6cedf81ad8228c0001},
  '{445, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'h00000000208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 384'h6bf105611bed561bd2f71d1ef2d6163a1a61965aaf7fe0220077ba91ac41c4f437bbf34135f78f0d6c9748c8852cdebe, 384'hed574398675aca014863cacfc6d4829a0f3adf8ed0a07ba7830e5b74c3efebb595d5f341a917562aaa6f76baa232014a},
  '{446, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'h00000000208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 384'h5c79378ac41d75a8799f8e2f41d9734ff5a3d4c2cbe0531d1e4da86b23d28add9edd6754b920514e10c1d3e091a876e2, 384'h5725b3c6ae8a001fe23f6f902df8ff5ae3721c5b790d7a61ec893df7dddee36fcc09eb01b19b62bd2dd8e1e99f0902f5},
  '{447, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'h00000000208b3f5ad3b3937acc9d606cc5ececab4a701f75ed42957ea4d7858d33f5c26c6ae20a9cccda56996700d6b4, 384'hea45d18c2d84646ad4bf834ba484909e79d12a8acaa2e218fbf81ef662ad3f3ee5f044dea80f06f0fca384fcbf42f208, 384'h699ad37f223aba03daf88e1a8bde46a871231cf56959d23760baf0f363fc8de77cee6909091c58a7cba9419d50928f94},
  '{448, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'hffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 384'h82526fe3465a1a3514c0dc39fca27eb0fc2c7a8666f8dfffcfd1f809d621f3bb775f2df3fbd9434bb6b99e1693f5037c, 384'heec53fc8b529a4b283137e7136317d77577e942f325fe1848756818637289bceef76b699b7eee6181b258810f910ab67},
  '{449, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'hffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 384'h33f8ce53cb494e377fb351edd3a90e6d8a82007a39686042c35137e5f6c6b50e92ea6426dc07257f4e2833669c98af50, 384'h9d3c8aea4d601702791480fcf0c9e28e757b0457bf64e9529cef0a29f2c4074d3e7b2d838ecd311334ca671e542c841a},
  '{450, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 384'hfb01baad5f0b8f79b9cd104d12aab9310146add7d6b4c022d87ae6711178b94d618ca7b3af13854b1c588879e877b336, 384'hffffffffdf74c0a52c4c6c8533629f933a131354b58fe08a12bd6a815b287a71cc0a3d92951df5633325a96798ff294b, 384'h38897bbcf7f806e2c7d32d9376462b0ac097717b984b3acfdb66cba4d20f2ea36f728342c21e6e9aaa517416c2ded860, 384'h0790f3b0f4a0c567ac9f58fdb42d1fc77ec08fc347736661cd73dd37993baad45af89a26d4154a6fafd81b4bae060e92}
};
localparam int test_vectors_secp384r1_sha3512_NUM = $size(test_vectors_secp384r1_sha3512);
`endif // WYCHERPROOF_SECP384R1_SHA3512_SV
