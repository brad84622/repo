`ifndef WYCHERPROOF_SECP224R1_SHA3224_SV
`define WYCHERPROOF_SECP224R1_SHA3224_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224r1_sha3224;

localparam int TEST_VECTORS_SECP224R1_SHA3224_NUM = 60;

ecdsa_vector_secp224r1_sha3224 test_vectors_secp224r1_sha3224 [] = '{
  '{144, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{233, 1'b1, 224'hb15b000000007c90bd7e479a53d6896b278efa828e9b33ef5404cf36, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6222915ddf6e69eaefce3ebda56ac501428b3d69b7b94c0e9ccf0010, 224'h5acbd1d130b50c08778175172a9d0d0e0e36b6a68c80af9aeae41b6f},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{234, 1'b1, 224'hc7e1590000000057642ff6b9373479cc4637154239c1863c1743792f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b8e3edaf6aa9e6322e916ba1cd2bce6ce694ca8e8f9f999efe9cc07, 224'h793b8d557b98e504bf05b2a57b1fd1eaffb38eda30db7c5e8a559c93},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{236, 1'b1, 224'ha84aefc841000000003361df1f290d1692220b091782a92e8a363329, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h33529fcafcd107596f846563605f0d9c479f5ac9498e325e034fd001, 224'h75e231e760bc10eb97901c2b8ccf908099ce7fc54472fcb419784d36},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{240, 1'b1, 224'h00999f1686b81b000000008f0eddfef71b4a955f469f2d3f9c601cae, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h09463baa1c7630494a9ed5d64fa2fac19ac452b3142f8bf19f585574, 224'h3897d58b8aff942a074a583604b174ddeaf230d7cead58e74835d89d},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{241, 1'b1, 224'h229edc99f5336a9b00000000d30aa317135d789ab8d4bc7001cfbfd2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4c2ba44adbb44f6b0f57de21830870d5acfc68e03c8f35e1dda14cec, 224'h6aff00cd6417ac43c1ea7e107fcfada404b88f4a79a0d12df96ab028},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{245, 1'b1, 224'hdafee08df93849e39d8f36a00000000055074d4f2f50cc395cdfbe7d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4e0f67b081cd6b87e3f4d792f1ccdd66e780d8028eaeb5c40047b615, 224'h14c42ea50c712c3fb7a0e18fe06b23822e9063f15bf2759dfc70383e},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{248, 1'b1, 224'h533901ad04964be8aa1f86740c274000000000c3445bf8cbae9dbe88, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h11974f58c95f8c44522f8359ae5e942577b8fb575a2ba18ff383df71, 224'h6c141327f9e405729c300f16b301de140c8df92c05637db952216e4c},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{254, 1'b1, 224'h32206da1548d2c97eec2755f5fd49ea5e76a27d61c00000000086b63, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h023a1d2a8e49deac352acb3a6a758070b5c8a4e75fcbaffd9f32e862, 224'h5d2d511ed37cf7d023a5335c48fc2f63cf0733a1a786c49ae929ce5b},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{256, 1'b1, 224'hb1590f4891953a511c5414d74383e2e54d811a36d25f1c0000000040, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5c845a275521649bde9e3bfa07d6ca528f6e143d19e97b1e9e305e71, 224'h60b4bd522c44b4c32e87b11b6b80b2061da98b4cf5c56dbf5f0651dc},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{257, 1'b1, 224'h7f3932b8f1469bac9ad91834d5d7f1f792c68187adf1fc6000000000, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h260418182c819de5bdb8851c5ac937ab8d83ab70640010f7eeae13f4, 224'h034c2f5ffaa2b4f1f111f4758e5adfbab5b7cfecfa48c8d88f5b6816},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{258, 1'b1, 224'hffffffffd9f963c65ba7c514c1e5181bcdb839ad0cba69da5d60a561, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0346d6521c74bfb34342c4b03c067d3cdfe35d3ea121580668301431, 224'h571dc84cc071e25b98d47c87edd3f6db73f995e5a4fa038760c43cc3},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{261, 1'b1, 224'h1c7effffffffe6d0757846274f00c3241e3dcb8e50cf2e0f30f36fc4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h43236a22ba681bd71f99a8ee2b425b784ba6ff55cae154bf1b8ef454, 224'h09cffb77306a5ea7675578bcfa2d2142c9dbd84401e09f78ec29fa74},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{281, 1'b1, 224'hb6951fb6ca933c00668c1b58f396987a172ac34bf9ffffffffe58278, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0c6822e256d0190b4962c5b4bfdabce10d277cd347caf0850892288f, 224'h3f59727e4d9e3b92f4b0ce710c5112caa18e4051cc71450f6989cb9a},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{288, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00c359b31b3ee10cc0bab7d21f0cc5cecb632186e8ca608a74f921986f, 224'h27787cc204c5ed561897c14961f7827b5f97395996de6cff87862771, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{290, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00fc0341bdbbce3beee1be9f02e46148af9da53128e0e3c45af1abe4c7, 232'h0092acfd718352e7107fe08ea6a35d8badcf54f57065dc4e8c9f2705d2, 8'h03, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{291, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h50b14256f6ea50d9843bd9e2b4c2d9daf75f76ac4e4e757c712b3053, 224'h594d68e1683ec977b2efcc8a7ba6c46a0e6a668a03f4f50a3e21e4ce, 8'h03, 8'h03},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{292, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h7801e48011fce2685a2f563faab34fff728ebb6e92eb029fef124eb5, 232'h00a9be2c1b86e99e44ef60e6c02a04a16cbd968482ed2ec4c1463efeef, 8'h03, 8'h04},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{296, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00ddf53cec8d9c6062904d2a04f790f4596c67696dd4f5422a3cb84c9c, 232'h00af10f2d1eb0e0ff28fa8e40a91d8d4addb20c085d635158de1a67bdd, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=56b(7B), s=224b(28B)
  '{297, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00f43b4a87dc12c65bf27f4b8610486402327adc0133c1db8adf4e3f9b, 232'h00a61aadb4c58ac0b5518d1c2929068eaa0d6a5d5f84dacf66e5b276ff, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{301, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00af736667b618cfa5526f073f7048d5e6b672a05569cd2912bce8914d, 224'h6a030aa73fd79517ee8175800484f2dcebf02871825cc67c41b1a8fc, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{302, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00af736667b618cfa5526f073f7048d5e6b672a05569cd2912bce8914d, 224'h6a030aa73fd79517ee8175800484f2dcebf02871825cc67c41b1a8fc, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{303, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00aa2f981add5480e7f2a8ae50fc52258612ad6420a1a2cc2c252c1693, 224'h32c1ff19c331d3e52a98add7e7f4f8ac122ca961b8cbe4260ed83e4c, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{304, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h008feb4b153b7dfe4081069ec708fdb161716ec3ed17c81efb1bb3e396, 232'h00bbc90cfae2c3957f2cec75239445239a1c0e9e0a032385d063f1d2ff, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{305, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00af2a29d356133f4d726c64e8ff7d80851649cf3e35d2b9de2725bbab, 224'h6d2199d9f3e0f0863e671deb987afdb25b6e6b7744bc53faa15cac53, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{306, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h7bb0bc9529b06a424e8efbaafdec5aa339de5599f82ec9e195f0cede, 224'h381dc950caa8b0454fab70c57e06a15bc771b693ebb4013bc85b56ac, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{308, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00ffd40a19c09ce0a21124f163c72558e1f15a11aecde9dde08c465bce, 232'h00e3cc54426c7850ae17670e1cc19931e9d934610f42f456b8472a8047, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{310, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00f480a474e28f987e1e76e73c7a9c5c12307f5bdc99d97e515e71ae42, 224'h0e310ab3403eb44f8f17e217914d136c8e2341f71177052d4f07dcb3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h04d2a54e9e42beab49a152ec0764b823bd92a0bf4d6767e261bb4e3d},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{313, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h009a24375b03b78c20230867b842c680bdb88604fa93f7c59317348310, 224'h60090ff5dec7b6fb6df459befdfc5e9d440198e8610a267daa9548fa, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h79823515d525dc02f18810142537553a6da56048fb999d3fdff85f70},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{314, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h71f01e6070a5bd694092417f75b1f1b35457421e9997fa5086dfef4b, 224'h2b8f67510ac820380907503b3bcdb89fdb5f2688434dba79d3a40a11, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h23515d525dc02f18810142537c3fc1ffd9a43852c262974a2a1640c8},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h453355214278474735b32b1d45c9a203421578c10acd426e9a569d5f, 224'h6b5655138346d0bef9cde0ebb97b4938e3c28dc612b4eaaba862182d, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h46a2baa4bb805e31020284a6f87f83ffb34870a584c52e94542c8190},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{317, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h6fc6ce348cb17cf57fe18e21ed13e8f33e5a724bf87f151ea7579633, 232'h00bdd1fb53ba4ec9a477a6f3e5193003aaf462c857bc4a20bb62446552, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7d96ad58b0dea0aa5b2f5689fc4d2f3f919327bf633ae0b17d506e00},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{319, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h3ccb08210d0b2283f3ccb779079bb160cee3cec9263d356565f770b3, 232'h009fb0edb83cae0b730fddd5c0d63e10a99e527497a58c18b84dae8e8e, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h78c4080a129be1ff118e039df4e8771bd400870015d378cf1b951fc3},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{320, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h2dd3cd29db7616a6dc77bb1a66e849133b1408c540ee2ebb01e07bc4, 232'h00d3e5786401c4533e15697c6bf86e14def5088590c19aec9d96f8538a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h5f3f6b9c25e45c8089f2c6543d345037e17f2f7d4b7854ab399ee32e},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{321, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h53e89d29406622bbaa1bcf7c980d523209646cc20a4b3104aa344264, 224'h7781d3de43413dfa061aa9b2d7c29eca9c8ed42b285fbcbbe016cc1e, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{323, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h4b1b3c491443d1a45cbe5fb2f6ed36ac3ebde2a2456a7f9afe628dd7, 232'h00d328db165ee1110765797569b30b041984790ea3aa65bd0ba3341818, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{325, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00d0c80d942da3dbe662467e1bcc69ceb322dc311152bf15557ed3f7af, 232'h00f7b627b0ba59524170527cc1161abdfa4a4a25dfd09c59a98db7ea04, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{327, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00931606b9f180d16409efebc996bb1df442b84e19bcc9bed0e236cb64, 224'h50edd2162625a979a25b231fba17878b756a77c167223886613afb03, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{329, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h008a46670a9c9d3cf03a9e9d48525c75e572680a26278adc0888d5030f, 232'h008c88e59829d5a802c0245aa8b5641779877c5647ad2b9b2a736535eb, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{330, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h16428097e6eb65688905678aae661f3d83b7e5ecc7787ed22fc029e8, 224'h68d62cb89be54d10ca5b575aa86f9c8fb475c6d90f59d4477595c01c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{334, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 216'h25094ea9e4ce76d8c47356e4ae604eb6469669b0161fff805a765f, 224'h6f807430f186ba63ffa0f315be721ec43baef24b8fba10b04f19189f, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=224b(28B), x=216b(27B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{335, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h754267d9f090524d4c97bb1a5622e0c9f804dfd70cc68d9872f0a4f8, 224'h708c24a49b81307db458c020fc7374770858faaea1d6ee37bf7beae3, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{337, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00d357674da166e0f4a058203df23b8f8ada82858034355d23aff5a812, 232'h00edf6d5265ed40b6da2adbe9f8cb6050ebf61ebc0e56a10a1d6cf6e2e, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{339, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00c1678bddce5f00e4f41ebcab86f801b4dc050a1b2da8f9747b5abfc9, 232'h00f1cf0d67d9c93456988a004dbcb8e95d17dde4070577e51d881d8859, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h09d2cfd575986bfe1a7420c7dabc0476e0dd13e54e01aa6f97b9e027, 224'h464ba5b84c4d92ed9fddd0bbcb2382f0e9b9d5bb201b2ea8eb8d3a50, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{347, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{349, 1'b0, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h0e77efebdac83c01dce3f8c4162e286b38b7e23de83637a72531eab7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{351, 1'b1, 224'h6b4e03423667dbb73b6e15454f0eb1abd4597f9a1b078e3f5b5a6bc7, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h474b086cf4754c270d20f88be569b7d7b6eb6e55de6ce21382160e81, 224'h60692fdb35b4cb824a2729fb175f709d06bc9f4e8bbb4b1058c53788},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{354, 1'b1, 224'h9629e241405210082c4e5e4b5925464253bec320eafa95b4bc5e40ff, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h6efa32457e09b8abe22168501bc4ae051d2294674114a9dca94c51ae, 224'h3173b652c78324b877dc5bdfe80324aeb01b171fd2626124a44f0b36},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{356, 1'b1, 224'h5d7d45b46692e51f9e2bb3f3e9f02672c85dda1d6aad741de70b0255, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h6f138512bf05addbb536b976b9125e1228f43f32f766325d1c270e16, 224'h556205464ff65c9a5d4d9475167059863835644b06862f1b49cca20c},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{372, 1'b1, 224'h5d7d45b46692e51f9e2bb3f3e9f02672c85dda1d6aad741de70b0255, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h3186a92aa760960996aea13f3137acf00b82b2b2036e607ec9c44b67, 224'h1835944e96b6ca1f445cf3350f105a97a37252f85cf6d8e628c96a02},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{380, 1'b1, 224'h5d7d45b46692e51f9e2bb3f3e9f02672c85dda1d6aad741de70b0255, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h500c9d08a0ab52d35fe5cf9d4eddea0eb8cc00e8e8db0a29a512de10, 224'h482d0f78f2808e83f10bee9fad61f4bdba83ab9a4f7d71c9b7083e13}  // lens: hash=224b(28B), x=232b(29B), y=192b(24B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224R1_SHA3224_SV
