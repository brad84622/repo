`ifndef WYCHERPROOF_SECP256R1_SHA3512_SV
`define WYCHERPROOF_SECP256R1_SHA3512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp256r1_sha3512;

localparam int TEST_VECTORS_SECP256R1_SHA3512_NUM = 329;

ecdsa_vector_secp256r1_sha3512 test_vectors_secp256r1_sha3512 [] = '{
  '{1, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 256'h1202069b6b5ffadede2fdc290da1badc989ba98a9a491db339bfe478450ef9cc},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{2, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{3, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 256'hedfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{4, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{94, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 280'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d0000, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=280b(35B), s=264b(33B)
  '{95, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 280'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b850000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=280b(35B)
  '{99, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 280'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d0500, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=280b(35B), s=264b(33B)
  '{100, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 280'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b850500},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=280b(35B)
  '{115, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 0, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=0b(0B), s=264b(33B)
  '{116, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=0b(0B)
  '{119, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h02dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{120, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h02edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{121, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57efad, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{122, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b05},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{123, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{124, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 256'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{125, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 272'hff00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=272b(34B), s=264b(33B)
  '{126, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 272'hff00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=272b(34B)
  '{129, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{130, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{131, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h01dcbe02d28091fccca712175e1effda760d08c16699295b22355e5e3ae9bb147e, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{132, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'hdcbe02d48091fccaa712175e1effda76933acc0b4afa1e184deac8b4f0f4c9dc, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{133, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'hff2341fd2c7f6e033458ede8a1e1002589afde39470dee4362be5b6c8812a810d3, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{134, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2341fd2b7f6e033558ede8a1e10025896cc533f4b505e1e7b215374b0f0b3624, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{135, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'hfe2341fd2d7f6e033358ede8a1e1002589f2f73e9966d6a4ddcaa1a1c51644eb82, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{136, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h01dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{137, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2341fd2c7f6e033458ede8a1e1002589afde39470dee4362be5b6c8812a810d3, 264'h00edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{138, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h01edfdf96294a0052321d023d6f25e4522e1324bd0b3e61f56adb3b10db3b750d6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{139, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 256'hedfdf96494a0052121d023d6f25e45236764567565b6e24cc6401b87baf10634},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{140, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'hff1202069c6b5ffaddde2fdc290da1badcdbb4aedcf3317f2e460619b548abd47b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{141, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'hfe1202069d6b5ffadcde2fdc290da1badd1ecdb42f4c19e0a9524c4ef24c48af2a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{142, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 264'h01edfdf96394a0052221d023d6f25e4523244b51230cce80d1b9f9e64ab7542b85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{143, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dcbe02d38091fccba712175e1effda765021c6b8f211bc9d41a49377ed57ef2d, 256'h1202069c6b5ffaddde2fdc290da1badcdbb4aedcf3317f2e460619b548abd47b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{144, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{148, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{149, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{150, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{151, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h00, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{154, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{158, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{159, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{160, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{161, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'h01, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{164, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{168, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{169, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{170, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{171, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 8'hff, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{174, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{175, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{176, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{177, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{178, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{179, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{180, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{181, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{184, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{185, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{186, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{187, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{188, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{189, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{190, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{191, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{194, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{195, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{196, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{197, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{198, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{199, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{200, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{201, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{204, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{205, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{206, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{207, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{208, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{209, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{210, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{211, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{214, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{215, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{216, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 8'hff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{217, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632551},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{218, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632550},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{219, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632552},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{220, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000001000000000000000000000000ffffffffffffffffffffffff},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{221, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000, 264'h00ffffffff00000001000000000000000000000001000000000000000000000000},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{230, 1'b1, 512'h940016e8f13841a9f29c65adbe20d7c6ac3d2a8817aa34e44be00ccc67db4f935bab243b106b6f3d68b875b328a96379ad7491c16643ef7d37225aaabc79bfb8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h64a1aab5000d0e804f3e2fc02bdee9be8ff312334e2ba16d11547c97711c898e, 256'h3d4e6c69176bb9e30eec304a30d982cb3f6073a2273f36b67b1b284899b08163},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{231, 1'b1, 512'h0000000097ae34ada66084471ced074cb11f6012595501e4f88b5ab4526808fbaabfff3975c6cf53455cee950965a5b5b71310c8a1822cb5d15b513b43dc5720, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00f521807c1e329ac6df4df24208d1e7088b4e4de5a82ed37dbfd8d49c7406f91b, 264'h00c44f723038deea858a25d7264d1680b416ffc0d909b94def9fbda02477d69ef4},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{232, 1'b1, 512'h4a00000000d34b9c928306129f1a8059b199049f30ffd4d5b9747c848b197497634fb5190298af2f6a90d273164d68431c984e0fcd3a810ccd7b95b5e0dcd21f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h219f842783028cab66f419241dee39da459e2d295d0ab1e56b29b38f50a8bd51, 264'h00f6f357077677e2669c1e289f65c6094c68b8e1efbe4c87468327c81d55979bd9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{233, 1'b1, 512'hf25200000000600b35bfa47958845baa9428119e3a1641db59a3b72db0b47470dc44921ca1826d81bc2e78142986441cb6a6c15880383e1ed77282f966ad17de, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h15768c2623e7093c7dcb468d430007fc7338f1cfd058fe22ab09a451b61ec34c, 264'h00a609689226f073c968fc46336cfd116edb92045f2383d5376ff88272dc444ca2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{234, 1'b1, 512'h9e93cb0000000075ad177fa53827e2d0b2d93ab1e6b099c341864034009c13d5ae494352e6106d44bfde1e40f82fe0bc542154fd54365234bd13e0a0e4cbbf31, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00bb449ace6f3b900103a09357cda16e3b14e9e99beb3b8f1928f0a66ce30b0ea5, 256'h6e6b65f9798cd8c32d7068270800da5d98f06d36836ccb7c30551717fae3052f},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{235, 1'b1, 512'h6d22e20c000000000726c9469eebfd2e764c9b4750557869e51bef687b0b07862ad496e4c6a056d46f5d244f5f10ad0005ded39047ab8247ec969c4e42ec2219, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h589e10e34c3fea59478a9301bde976cbd56ac15afa2f13f14f310e5e8d6bf1e1, 264'h00adf5198111939bd395bd3820742a68ae97f8595cfc8b7e1892fc360d13142158},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{236, 1'b1, 512'h5a5af3265a0000000025640fd363bfd88cc171f1966b1906138185d763f0ee7065ebd2a5813b79d02ca118763c60dcbda580f5ec322cdfb2c0a407e223f6b16d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ad5a1daab3023a651b58e3a13ebfaefc14fb9c79ad2610be68e49bd3992e5722, 264'h00cfb91fa16a32c8724cef5714e72f2c91b1d50050b4eb272a82327604486cbbb2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{237, 1'b1, 512'h6c0f86f08b1e0000000069a0652407ab389f7f275bee385294bfc2a7a9119905f5ce4e1af41b3850d665c942f16914cf903717ff47c4e186c7fc97496a068b91, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h59d0df1176b277e12c097e9e00860dc4ad3bb7f2e4af2282beb13eff9d7b6afc, 264'h00d3da4f61e8adc8449885a52bf73eda66ac1b77ba05a1ab8397e42ecaeaff68cf},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{238, 1'b1, 512'h5ab9d448ee67ff00000000baa93e38832a2709f7238f9bceb67b53fea917f665de9153c44b7280e1a5674dee745f5350bb3f2259ea084b398cff74d33bded951, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00d274baceefc72a921fc4962cc9487263ec6984f0f82c0b992ae3c80ba685b423, 256'h24bd9a9f39ed02773e8ba54e3f0f99f4e806a69839b7890099be2978cd55076f},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{239, 1'b1, 512'ha1eaba175145939e000000007804c10bafa1416c6dc9d3311f844fe42868c6bdf283b946814df78822f198d26d886ed4713421a20dddcd82a21333d922eb39a2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3411db9e53af62472c8afa3a4ae7d044fdbb78b1e3a8e8fd329bc72e9e1dfb5d, 264'h008284d93b62242f6274a26a3419719dc0635e0604fa6da5c2dbfbb85541c88566},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{240, 1'b1, 512'hb1fe8fe86f9994808c00000000f313a999ae7b5281bcacf933f05e4c8d526e761afa3141e9efefe959438620220c28bbad7047a6c1a98f95520baeb1d7af6278, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h33b2abf92021a14fd1e5293008c8aff551fd4a0cacaf8ec6e147f40d0f521cb0, 256'h4d0d3ed085477a4dc7fd86d242905637a71700ffd4c22cf962a67e9ae32b8877},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{241, 1'b1, 512'hfa3ef856182ec646db7300000000241a0e98fb88ce661de43bfd86f1c929391ee9ce6c05612b1609d6b8466a9c4d0af24ccb440f463cd18addf4674adb2f94ea, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h717f5185242ac57215d8713f902cf9012f45dba76b8e7e51c67b71e6de10f0d8, 256'h28a9ad765a6b1248807be126b9eee01e8e2d65d8528cb28f0d45763f507d97f0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{242, 1'b1, 512'hed19e69c6f4de76b35ce6c00000000ad94175b8ad5f1fb69995d7d87abd893772b81ff83fd6caa25d1fe69b0317ec4068cdddac49512e6bf12d9cd8ce9a951c7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4e57dbece14d3d279f1e831777b28401d2990c4ae477eebb997b583e82f29c54, 256'h3e41fe090c8f14b8af7fd39c2628869258cf05b0e289b6692602c10cdcc8dd83},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{243, 1'b1, 512'h2e2e984df4c5b45f7e337184000000000600f130d66940e8b4c0c1030e71fb8df7efce69100b9174baac3e7c474054e875f26cc182e925a17f55688964033e9b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h09eb0b2bf6a2491eb35c3a902da3c6c90933dd374dfb1f60f8ef7bd749725755, 264'h00df8a0ee8f757dc599350bb0e2aec515451152ff05bb2e439ba9145fc9a0849fa},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{244, 1'b1, 512'ha8f658c6632e4f474a6f1af1b9000000000048ac2a6121c8add714fb8cce854dbf1871b07a75008a42baa6cef01b4875eba4bc9327b41503cb36ac20f9354238, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1c66a303f7f548ff4c17ce6c6038879cb9d47abbb71ad69a798d0d8a99518dcd, 256'h485ee205c6fa3ffe5411948dff2351ab9bbbc20ca419d6182da77f5579058749},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{245, 1'b1, 512'he89af705f005a4e1c5983824150000000094795c26507ca965c1eaf5782dd829a5fb5464eae46688a19ca7fe5851291f76fcd7f7226131d74cb4dde6063215e8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ae1fd2dbad7ebc2b7f19d1789e1f68ce345f40568a576a29dadcf894c51f7a3f, 256'h69e80f80c76b57e1767484485915980b5e2493e89d8824b7922ea2cbc687d2b3},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{246, 1'b1, 512'h9490ebaece67e31eca85b20871120000000077b2785e29958e0ab90faf8fcca953b142d51892ae5362246dc07a066ff6a4c9fed90a79fb59abdb7c8a888a9652, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h67afdc527b0003c8400ade54df5663635f811950cb34ea77435c0ce400365249, 256'h7afa3d39b8a7e52ce768e466db6da41a354c12ea2f677bf05a24fc689e347323},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{247, 1'b1, 512'hdf22c290212fe9b66a9c65575e7be8000000002b9d4a3251cc7b64eeee3e76b7e65ac253a2e3d18658634eacb7494688a1616feaa0bf8a6cc0edbdeaa4533490, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h009b1a90f8116d33d674137579528f395ed13ecbc238940a1a9a8504a72568a9d7, 256'h07f34d9400af004fd657144ce97a13b76d509f7fd4c9245ce54609f749ead3cd},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{248, 1'b1, 512'hca6a7cd52432b20d8cc73c4e810dc325000000006ee638ed6bda85ccdf3b4606a300f2439910d382aa47f8e5839698e4bfa1756c5e93b3d6aee97edbc8ae7794, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h263040f9babb63aec7d73fdbce988fb3ca2115ab24bba0c80832e3de34b698b9, 264'h00f7d99b7738aca745b91b65c697a83ac76ce1e61568d9271631d06af1b77ad5d6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{249, 1'b1, 512'hd912418a7d72e83ab66eed185bd627c70b00000000a88db442365b3ec21269abd09b4b2e040304518850835236add11fecca5a2c529f8bc4c06174a03b997830, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h0082f676de71ecae7041b8788e0870a57923c71fd21db1f8864e4519ee2f65d888, 256'h020f12d98b79d45348513696d5b4926856d953e72f267d30e7bcd57ee8147210},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{250, 1'b1, 512'hd8cdcf759b329e28b173d8582d7a91bb2d12000000001faab0678de44c1caaf5247d111c9e465596a89073d5492cadb0bc766620952c817f31a391f32fb27346, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4e3c9c22a54f1ceb9336b656bf7019c375cb7f9137d692454c6d882927f16795, 264'h00b3bde8f45d5f885948b45402b9e7a722c292e88bfadb5bb2fdadfe8e1b3f5181},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{251, 1'b1, 512'h91f07f1a3d4b600628f1754ae5ec28d43554a40000000051e8c4594c5a2e68bf2f497bfbc7e703e1b18398a0b5515a38d60284b1a2dfad8c9132a7b9a98db6eb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b20721bd0e8c9ee6eb790cee9d88481d17d568b4c942ba437e607460031c1df5, 264'h009f13ff6a54e6a0c5041cc3690c8f3b499f05e34f235c8adf8fd455df4a17ce97},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{252, 1'b1, 512'hc6208a5a5c6b71a957477d8c39b01e072a65ac1b000000005c6ec3ddb8ce20911bba1864112d3407082c700820f8676037efb40be95619c9f686163a4d0cdc5e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6b1d46eeacccf7066a0fef27f498a59a9376b2544258510452787bd4a35783b5, 264'h0088328ac07938b5b9cfe62a3841382cfbe9d623480cec2a3fdb73ee36dd4aef8f},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{253, 1'b1, 512'h7da7793b2bed3ce23ef7f1c04376791fa03f741f650000000008744fe10ac37fab4edf76492a339fe79e56ef75aee6c3169a0a61e3cb27e74666a4fe4184526c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h257e760a54637387b443f829f1a5802c7fc92bdf033039acf68e1acea0cbcdbe, 256'h25087f120467a80cc07efb7bb27ae68d8569a38fe2908282c3c7a310322761c5},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{254, 1'b1, 512'h48cd33f55583315ab2131d5db1f9cfcb0590b13a266700000000c9bd5d6fbcdf457e3bffd7b4875145a47be68b99a201b93b8685e80d61ce692a913be1183569, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1869c821e271838453c88c4a867df2301d27662b72d9385bacb6740ab6d6b5c3, 256'h22ccc9a0493116556d9ffc7582253c581452d717a7e00618dce21f46f5b64fd0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{255, 1'b1, 512'h1acaa001f6ed1b1a5b0bbde85513fe0b7aed266bd9da3100000000dc1113ab87ae3bf815157a1926b7bc3f659934702113570c26bf1bcdf1c8492f79614e844c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h0094a521fb3bed347b0dcbe55f2e67c0d7abc4aa32ed2e1a6fd1c209de3a25ca25, 264'h009b7631a6520ed4b14b5b2a8b57a52de31f583b8d1260eb8dc061ad965d0e9eb6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{256, 1'b1, 512'hc6244ad67598a847488d31d513fc9dbd21d96307c296a4170000000012f527d2192eacdb6045c48c250e317b7fc62ea79321783ae0f400ea4a60b48c2a2fc495, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ee4913a5f83dd3310e91595ef197075600ae17785e1c0b9139cbaea8def1d6d0, 256'h2818f7847c48a9a38739c71653919104db8920a816000ed21e5179980efb6b6d},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{257, 1'b1, 512'h90f9b7739bb1699b90bfdf7cef079649e3f08242a08d05026100000000d3a4568eccd5ef4d94de4885986b68670617f552b9cb2a6eed337392b49ad4d04a9dad, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00e912b0e5436db2a50817c6424291ffdd41352916e956ccad9068c95125f3a1e9, 256'h73309aa384c56486b6a4c699fca446e6f67a1133892971be83b4e2dab49afc2a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{258, 1'b1, 512'ha7ee711aed6f375a8a15680f30deb6946501624b70b47c79d5a500000000ee6f7f0f2b69cde1a389e3abe86e51efe844c8e4ee7c3b2a15925d8c9b8b296ccc53, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00eb0b719879b2fd1676b3f6f913e353c2b4dd8201facb067e15da1dae9addcc8c, 264'h00a73b3a703857aa8d12263290366a19d64e0b3efccd0623f53a7370099e9dcece},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{259, 1'b1, 512'h9583a32b620d5614a1c36e06ee45750fd69ef561faeecded2ff5b4000000007bb68b2b419fd574ffe1760fa0203fb1718c4e5d8a798563fdd98439f37a56dab7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h0095617b71dc18a99e96a95ab5384324bff797ad704dfb1e2d6b3cc06e76652ced, 264'h00b11bc49444a2e2635d4d9b1bdedeb61593b5f3e0e16ce78da813ff64b728f8d2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{260, 1'b1, 512'hb6e404060dcf7182366941e77a0f0b43737232bbf9f73865863c271800000000a4ea51e31a92eede7497562eb5eff19b08310fdcd46cf3c22e069110aedc21a2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h28fbebb0c142c6d200bfb173173c03bc3aa55da6d48c1b784628f2b9f59038f2, 264'h00c0f1427005a46aac00a0af43b8f54a951e673e0480c6bf7a6b5775d4a3de5e60},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{261, 1'b1, 512'h57003aeb6ad8b84b54cdddb9243c65d8fd07ad1ffdd35f11c319f06394000000000aa9393490e8dcaf1c1e53ab5a7b2dfc0bd1dff4d0fc1e0c9dd5cbb035748e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h457ff86369e4efd69592b161aea2b09153f37cf69006907a7558998ab34b38a4, 256'h12692ffc569849dc8e3b9fd2cd7c6f42207bb4c07832d490c9d35a702665ce58},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{262, 1'b1, 512'hb47f61cf42394fa1c4c8cea80b83e366e30a938140f793851af87bd3782900000000d7a39fae605c98c96e0a5b0e8a58e47c3b50d4905171c884a64239fdd901, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ac70036f6058fd1eb40dc6f58dd68ab56e73dc6841eaa45a83813b6aaf75fae2, 264'h00f70f7f0563c46a07d248e80a65f38532d5759f49fc104184fa6718ca55274372},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{263, 1'b1, 512'hdfe80a6b887fa09cbdc8bb94300a4ad38f0380331a18c0a0b62708e590dd3800000000d364091041bb72f35391e792802f5c23fd676d0775e56ac2e41880d92d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h59baaba3992dab0b594a2e9fbc4c344cfdabe7868e4e77f47a310d94916d30ce, 256'h20b16c383085ee74402157d4f2da5f7e3e995dbbf53ee50985d4f7096882edda},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{264, 1'b1, 512'h16d0d407630fbd8dd9af18abdbdb902051c86b156254ecde6a5f0a5a1510f99400000000c202a44b1c172e1436f2252d80f9ab44794b22086f877c3bd4aa5fb3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00aa567a710f7010718b1e02792bc63f9049c02f798bb319214c97bc734e54d115, 264'h00ddb7c78b45c4221db6f26e845f8c30be61c29bcf38e38abaf7cbd03e5af914f7},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{265, 1'b1, 512'h519e4709f22b7ec44e321f4d403bdde7f532392786df003ecda243880f79f899f7000000000e3e6d749c0a602d959e0fd13a8a491554d233b9dcce6cac4ff3fa, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h6ac18c06081a51ac5fb6d0a0735af510dd0ad529206e7fc0c1b6d0ea36cec4a8, 256'h64d49524cc26ef8eda21ad5f2c371203d6eef8ddfa5da7a6c37d86f29efc1fca},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{266, 1'b1, 512'h00ac9e66bf4db08b47a08e0b34e95e7ec2da8a82091479dabd2d57199b450dda70f8000000005b979f8077a5a74eaafe42ec70504f2bf8cd07aa23ef52c0321d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00cf59dfd67512e2d173a398cb648805fb41e3099f27a7867aa2dda50dcf2e1f86, 264'h00bd528be771fa1e52cab6d7485c5887befb378ceaf565aca0f32d2831a466959e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{267, 1'b1, 512'h2cd7eb20ee13fc351891dc4acccbc978161cc1b1e0cb95127485ff132176a972377cdb00000000add5eee3b407ef394da0255f21b9b8ca144d7e76fb075c6bc1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h455f1c4406b598fc828ddb3bc77df7ad04baad399fb4975f542b19aeedfd5a11, 256'h4e0555d9bf4211d3ab173e2e6c7edb990867f8f982f6afc1b4b6732ee96a0af0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{268, 1'b1, 512'hca402f2de7f990c5e1deee30d418810cd3a8707888fa5d54d3a5a0b3bab20144dbf37f52000000002a1f22f563f07cc9d066dfa8881777cdaf8a1ae4d43d6341, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00e1dc7a439633b9bc91d37a954943bc94e5f56a0442a3528fba5c6070cf25e86f, 256'h0376b7ff7601978a47bbf7d11c6844520a442ceb167aec3a0ddf36e150a385c9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{269, 1'b1, 512'h4386a89b56a955feed663fb88786a1c3916e8c65775648439638f2278c7d32c6d67f942e7d00000000d3a5ae2110db187684130f7aed62cb05159f8bb6eb1b26, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00aeeeef010cf97f324e6f89f3163656305728a573b885c52ec5973eba863a08da, 264'h00904c25f931e78e2b59fa9a138cb80a5c22341601a18501d364af361d69cd0bb8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{270, 1'b1, 512'h9a76ece71e15ffca113598c14654fea437156151bf5c8d47e15a6279ff965eedbe79fd4437f300000000148cc8ba720cd12a6cafa72448ec2cd6ad2852b2f703, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0e3798e441e787dae4bf84e2748abce913f362d41d59a39d58d89c889e52229f, 264'h00e3a002023296fe6d9395fc92ba31dd35c5ada42e06db01466a24f087ae70cdb4},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{271, 1'b1, 512'h24abce8b935764d6a61bf597db6c773145d5992485866070fe22cd0f6f871d53e72f6abbcac6ee00000000840dc44c1955185bfcf393a1786b04625904f03e85, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h009bfe9e09c40fad40bb442eb045216c20dc1282d3cc4ba77fe2e3db92d312fd80, 264'h008a152afa2164548b6edfd6610046ee001fdfb06555677c98bc505b6aef297d15},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{272, 1'b1, 512'h3fa9e7c5fd635a7b587b56e19e8921e7cdc6d8f6b1ff03b579b907ccc2dba540c1782d5c35e3aeeb00000000a610ad03b540240313bbf54453b27d3794341d59, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1531f9b622d3172f72096b8afc7278eb7bee49b72e1b948e48cc1add8f01e365, 264'h00edc803cdb54bd4c54b87bc69a42df3dd11ab56bb13d8b5b78642ffa9ef88d31d},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{273, 1'b1, 512'h4025a46ad55fab109832d892d397d6e50c9c0aaf7136c275c259a6a61333a7e139b394a288148e32c200000000a3d26314f0694c5db5058ee34dfdd8fc2af9f2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7973333617680ff89798c6b64bb42f436be7771887c2d14a98dd3397e6896e0a, 256'h11b70b23a62fd9ce1b27c1b669c851187c09e9081f0aa6ae011411425f694929},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{274, 1'b1, 512'h1e2fbff1179de8374cc3b5f47b00ade36b6494b8941aa810476c8b40e3ad3d7f5f60d8ff0d13bdc7683d000000005b2a7c0d9bb60d8af2267c656e800069cee8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4fc40e0b3dd49c4f259c5ee2ff271b703b9b7380455167e11360bf336f72c0c4, 264'h00d219cdbfefa9ced843f947191ff11bfe4880702a4504f34b28481b424f433a38},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{275, 1'b1, 512'h1efc0d2c8682584f2504efc8fb5fd2848583ab11c97a1ad1d23db89d7d853316fd159eb4e2cee6ee4f2eae000000003ec9bbec801c26e55e61dbd6364bed8027, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00816c369e7b8672cce325dae1ad2f2a5330d177fe0da399c8e520f361ac770389, 264'h00858c9cdf1a2ca40ef9c1e02f883b34701dc1760a9d13ba714c57dd886282acd8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{276, 1'b1, 512'he68fbb72e90ec509836476f39f26d3f65c5deffafd5b86448457438ee0c621fc8f97e83c77ecd131ff1e33e6000000007c2a942574c7da923726d5304e0de79f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h51adf43cda1a938e1deb5fe08ab28df1e607f25fb2e98913d2579420b63056e6, 256'h3b8920181a8ab6f9ea0a1814171db3eb4ff3d5fd9cbd2d9c1ec4018a7625562e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{277, 1'b1, 512'h90bc23f7e48f29ee5cf5bda8b42a6a8aed3cb6018636758be3051cee87758ed5998aad924516e34c49319b58cf00000000b7f0c29548e1c1244f0caff38b285b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h42ce9e0f877b7586e7c0eb2fde6f7c4b1f4cc888f54402f2b7bb99dedc2b7f07, 264'h00f0413e7636cb6605e0d7284c7804d7c9a3cc0924d37fca7d4943d9e0c9817427},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{278, 1'b1, 512'h1c0e382d29f7ce824206c57f19794f9e8abe01e6af45a57dc9c01184c7b956aba27c6536c48c0951e2540bf566ac000000006db962ed4d45bf0d0c1c6c806b4c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4b2e5a797d240cd8c80b424a41dc47eaad249fc642e3c5b4bc68328fc1e26fc5, 256'h117910985597a6f7482bec7632e94676c432684f16f7f3d09a90ff4ed6ad36db},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{279, 1'b1, 512'h92cc3187d3326341d51f43165add210d496557c7a27669692c21c2912bc85d13d22a15ce9f2dc8052f89cdb3444fb400000000da250c8d1d81c198686e0c62d4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h42bf9a164723ef3f5cb59b528966ae648e80291785a4e0067283a7af59795bb7, 256'h017e1d24962a34d850d94187d269836ad437396a0ff134067b1baedef69b5951},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{280, 1'b1, 512'h0ec91d81506646053327c352b11803f36a38ba32d940cdec35246744477eb4c423fd81dfe4e728bea623290a65646d9200000000f68a3961185e3a1eb3a74496, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1ec06a62d69fca8d99473b8d5a8af3bbd701891df976e33e2f86c6084fb705f2, 264'h00b679eff436faa53c0a3c437717f574b59135d5dc49fb8524a365296db2d119e6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{281, 1'b1, 512'h290ba1c9dd4ce7537613a8092317a721e35cf33f17d8c82bc20a765683871857d7a7f0f72e659928158b11760b339f16fa0000000065c91469026a04f6e368f6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h183c81ab34a7d7c6742ede4198f5c75ed7fb79e8315899ef0dd26f95e3c4ba26, 256'h73f0196e459eb980b6e7ac44d868ab632d6421d1788b9f9651fb827b1a8e5dcc},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{282, 1'b1, 512'he9caa5454fd145db00275838ae34244a94ee61a025a174247c1b8056e6959c7f851f3038bc773457c88404c0dd497580644500000000719f683608f5718616e5, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00f5bec00e6b90ab2a8f188f8163dcdd9b8185a6bbbc623c12d583c9cf55c8e3ba, 256'h5dba085bd57b5471f8547cff0aca9e51234d85c0847d01a3aa0b3cf3cace82d9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{283, 1'b1, 512'h1827524c50d2a178cca81cdd33a0be182f764450e04af569ce80811e55ddf11bf9b04675631ccc24d816b26e407df93f288bae0000000040fb10fffd72f8f6b7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7c18891499af92cfa1db5538c7afbd44605b17dd0ede573206db85af23d3fe9d, 256'h28ceff96833996ebababef332b05372209844ddcc4c2134fd9311397e733b10a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{284, 1'b1, 512'ha5186acc06258c75ebd6c4985b00ae514a23405ece5e1c0a51122b5727c5b17a8adfca46c2479895b4121c304b5b2785c72c06a000000000ded1a008316d23dd, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4ed587536ba15e6707014f5ae773a423475e5e37564ffe91aec17722894cff34, 264'h009ff59fabe5e8dcf9539ea1bf9f4b880f112a26c915c14827dad9de6b251dd65e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{285, 1'b1, 512'haec77ef7d501e59ceb458f4b03194d730583d8282b6bb01ce0b0417143ca15c2059e8290afa26d6c1e38502d0b895bb4cb182dd4cb0000000097ca7caccc470f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4fb615772d56b6d1ba60f371eb04c557e0c9414c4eec00819c7647d91e7dee01, 256'h2623c6c4a3bffc596cb5f2f70a5a381942d350df04c35978f6607ddf7d57e4e3},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{286, 1'b1, 512'hfac59bb2cb17756c53956cbb809fb1dcf8f30340a8b21f7a25a1e6b500284c29820250c5c8492ecb2f1c5906b55dfabfb8c47b418d50000000000efa79a0e20a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00c53d6697f536b8fb0e79f3b002dc626a02948e206d96de7c62bd7f9736408ace, 264'h00c9423b8575e4afe16cfebefb03e55d628270264fad0eb67c9acf0268e514584c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{287, 1'b1, 512'he1942b44674c9c247d1f5857111e24baa87afe02ae74ac9d1ac122c10ced967b6243fd3055a4de1d50b98e24831c9f613d767a3060f7f600000000e5461279bb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h08012cfd3713068d8ba6f3fa453be9da95afa6572a893882075ed5d64d62a417, 256'h3c5d1bf341823a4cca251cd67d43a6bcd6b5e47303082b7e54c80df5acbbac82},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{288, 1'b1, 512'h9ea149f211e7bd1f624b20fd50fd2c474d627b16250fb6281c6bf57af0b868f48101c656162b5e1415c87cbb7a685fd752937f97cf58a424000000009deec0f0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008ad3da767111f41558fdc51723c649a87f58d42bea3431c8fdfa1f1096e3f2dd, 256'h7d1ea6859a0c932f2298f9d21c89ebea7354bbe508d2b73469dc3efe8613bc87},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{289, 1'b1, 512'he2d392cec1344167d947974fed90e637c5f80aba4fb00ba57dedea9f7ffd1b0404437d90e50f742cad5ed8b82bd136d13319934da1f04f50950000000059c93d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h62becf5afb08835f6768882c58a26c501f277ecd61a48d1fe683b6a78c49ce82, 264'h0089d11230de6953a1eeeb6b30774fc6bfd093c1e7c0422a7253428ba17ef969ce},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{290, 1'b1, 512'h40195fbc1bc4b600980e2c2b763857780d875bf68fa15558b038d9333a6c76f3aa4687e0325e29c3945bb8ac11ce675dff92bd5dcf0efe1264e900000000cdc7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h22b54382e2f2e6d7cffe3b34fbd567c8b503bfa6b5c3e5b8131e0ffe20747176, 264'h00a6d25ae5cab39cc83116d073cd1eb59d80ce2ed208c1c970b134be2ad29d6068},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{291, 1'b1, 512'hafc1cfa16e5549a03769a98e0a323b3ce3d8e3f316cd9f1007e4366b81a3affe3acb663d6a5d6a6857c736ce28eb85c432aad5ea98a80abb0b973c00000000b6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00e2d9f5c37ddb25978ed4727b63a5e17546292526877e903f11d3d29874e952c8, 256'h5c28ebafa2c2d285ed7f143d49b6d47daf12ad21c36f78ed7f18cb53d9c29f76},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{292, 1'b1, 512'he47ec71fc0cae21e08260f64fa9dc1a4c99ce92048144beeaf932a124c0f87a8b0db214e5424891f30a4cc0311efbb2d49807cc31733db9bd80f912800000000, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3b4c2fb773223c1dafa6d6de9ed2304dc25eea1fd487442a3a64ae8dc8f14927, 256'h56c21579e85fc9075c7601bd36ef8a3fa57d5bc7550c9a17bb8383e7fdbb366f},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{293, 1'b1, 512'hffffffff149aabbf287a78cde6477453f7f9c2310cd2d58ece43bb07019c69c965ca25e8df7696c97ee4ecd4966f7577eb41a60745d031a94f5856e1a5f95aa5, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h05276f6159e2853fc6884c2939997b5a3be7ae615dad7517d6006208111dd678, 256'h059ea3474bc6908c565dfb5bc72fd1a84231363cf78c4c317a061dbf1b03cc07},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{294, 1'b1, 512'hd5ffffffffa5bd8691d54adc06abeae7d4857cd52aa3ebae84fb391361d804a381d15d6fabbedebceef14c94b5bbcf1560bc8b97cd4c4accead9b453f6d27746, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5f856a30a8803a2276e8e5b8475f085d14f6de0c5f64eaf9e9b81c75fa831672, 264'h00a210a74c1c682de5708b9d19e6fd2f74ea047b1352edac7e4784cc008e8b0b5a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{295, 1'b1, 512'h9481ffffffff6e35dfab283e61e8f9a49de1cda44cdf1e2680292ded627b16d9b566ac057cef4c3380ee126c020a6ae86ded132faef613440c54185ed5986dcd, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h1c058daeb17f995cbaa4b02fc1ccf0a121fb7673d7b9b7bbaa2c9d850f9ba741, 256'h3e5400acc992698dbe9c41e25547c6ee08c841d6604de457558ee8af11d54446},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{296, 1'b1, 512'h2d8fbaffffffffb42e8498ddf2697ff4a2223fac0c486f05f57374d84dab9e8d13f52f6c898c8a7a74f2d48bee3cc16265e12a6dca3bee77c0ff0ee5e9af7e49, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7a6c6eb198bced25223fed630dbd2956c3799a21389e007efc23a0b3968f8aa5, 256'h4535354e8fb477d0be4a16f44719d94650ed4607eabe206848ba24322406c1d5},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{297, 1'b1, 512'hae17b907ffffffff72c833830a0827c91ae711b1704754016d3b0ef4c8367a7e93d4ba6f63e6bb8d572c24bfdc55da0d39f5fc8def9b04723ae25c1b82a3ed86, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h009d05a43f8dea2c4a3c0838e5987d899e63317a17fa5f609a4baa3764dac9899a, 264'h00d7c1833485f0a6914e5633115330a59b2ade5153b01b2a1af0a815f44d7f0aaa},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{298, 1'b1, 512'ha55ecf9029ffffffff0b0266df6f2fc70941d6389583046c5649a1740aae64600c31269408a3fe8dc0975b57d60cc95053b7d311b677bda6e8a0d6792e328bb8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b262a757ffcb496d880739d1937f139d39cde8e7ed29512a3be51ad470dcf5d9, 264'h00eb8dd006680530f27326f1c9c54e5c4300f1bca21bdb17245c485d7b296a2372},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{299, 1'b1, 512'h37837a8407b6fffffffffac5686980dc2ad1a556be4d1fcf5dc000a18139c2322fb6d35995be1b96f942fa8bcb31b6d4c0efcdb2febaad183b00f4967c63c04c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h480a6875b7bee4ed80f70206400df10264c38be42b07443c6ff19c0aab580444, 256'h78e3fa1c2fe11208c189a39e717b19a51f5172054891c083931861c7919d4745},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{300, 1'b1, 512'h148ae8a9d1f212ffffffff9007e49461386bac4123a9f847a6901d8d1508c822348ae29c100f38e169470e9a05b8cd6c780a06d49e062785dbdf1fd4cb89afbb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00f2be8cc615b14c289e50114ae2473b105447ec8c5311ecc3abcedcbeaeea1983, 256'h56ae20cd659370712e06bd6d5936bcaa06169737a062438c7e599bfff0099fb1},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{301, 1'b1, 512'hc17991fc38743c0bffffffff12be8c0818873e8d65ea350547aa4cdc067cd0a4c21e1d9387ca3c60306f95160cc1f85a08ebdd4f3107b359483b719f5b9a18ab, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00bed38f88fd52bf1cc4b4cc58bdd8a81af894c5a45bd822acf468eee08a683584, 256'h1c9f77ab2c821daa896e73b9f6ed4edf72ce62a6c48b5caae6a5ac9edd8d2953},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{302, 1'b1, 512'h45477dd24fb261b2dcffffffff376705fc972d1fc0eebc57960e96dbf0315340601ad9582193434f8cf1ff955cfa9a803a99d9465ab1d11337155273e65b2735, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008513ed012ea7a10d2239c209e172edb565b1bfd2cdfd80269f79956a4aab5af2, 264'h00a413070c1e974643e5d5fdc56209e1421a254f47fda3312ceda244064efe69ce},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{303, 1'b1, 512'he4d30dcc9e0b433fac32ffffffff83bb0169390c4443bfa7b7bc8a7c4421fb94a64d266b35ee622ee92a194a9c369a1bdd0961e4047a4fc3ed632b51f01547c1, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h25bc1c38b291a5f60b7b01eec8a5025c69723b183f9090150a7f0ac87464f2f5, 264'h00c986a03025cbf9bdfa4e9a0988822dae44c48624bc63a203072c9cb1b813102d},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{304, 1'b1, 512'h8f46b06e493783b6d3209bffffffff5f263101ceb63bd0313945c63e59a123011230ea2a874c147574859882f49e6fdc842cbd97843daff440629f6a58573ee8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00b721214cff1779b8f407f4b1b2b2c5aa4e49a4a517031ff3d24b5af589b28b96, 264'h00e9c53670e94337535dda10a599de0a6da240ea813e8081f9caa6bae59cbd310a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{305, 1'b1, 512'h34de554e38945bbfefa7cde3ffffffff7b63c616e7853caa71db174d8c61626ec0c2d1fc20cbd176f51bd580fb3d6dbee8b1319ce824b44fd820e94589a562ad, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008695064bbd15d76b698e4bb8c0183bc2634a5c2455d6bd2c3f8323a4268edfe0, 264'h00c706f66507b52d2c8865e3eb5959267307f51fdb0565c2320132f2ca14123452},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{306, 1'b1, 512'hc80ad608a993f311fc5d85b14cffffffff76d81aa75f097430416ac8d6d4e8f80858d995030cfd10467787a708fb59252ba27fd5cb768e2b3cf03a351aec1402, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00c91aad6b3c086073dafdb7688c6366be9127d9935cbc6e0c14b9f76c9d272c43, 256'h73c0f75156531aad36d2d14169c2b66797e8dd31d6f66b8ddb83f7522fba2176},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{307, 1'b1, 512'he9f4410a9857187394e0dbde1bc5ffffffff22ae4f317b16e8c82ca5e8ed1488b15705fcee61951d122b9603a8b3744eb429a850db99537b15bdee559ceb17b4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008125832edd19949328b170b1067eafcc17b3b79f5c139dfb6c109a1107ac76c8, 264'h00fce7f770e2245eeab16c33a230f6dea2ce1da67d11302a8ce7dc6145c30a2bf9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{308, 1'b1, 512'hdbab4c37e253fc1deaa9e71c035737ffffffff6e927ee1da438de0d1d5152cd6d0549d2b8172bfeb94749da7ff020aa760407bc5e12a5a099a45a301588b62c4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5e399962385aec963cb80dab6b5f5c341ce15e437142f4275ef9c210385348c1, 256'h18a8157a0976bb0e349a02134fad0d0286c40a5e43a47b49b5a03653e3ae9e19},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{309, 1'b1, 512'h2ad0f69e7f2e5efe8116b4b576a322e8ffffffffd986d354530161e2776001b50987f4eaccd1eaabb1c1d4d6c94e4f7460ebae1ff8cbf4a1df1cbf4a3e01348b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ada147d5937331d037083c0bcda59adb6125485a9ea78ef6884c1432e93e4093, 264'h00b5ea223b88f45533826a8b24fc91ed80ae3560543102fed1d82360372988dd74},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{310, 1'b1, 512'h69e08e9fa0546aec130be51f245d0daeddffffffffd8d24508cbc6106330bb7e4453fa88ddeeb7a8b80db338a7f66e078ffe0ee91d6b432c2d52b5a0a15f847a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ff56b22aca9206d8dba458507804c9f80b94e75d2b61443a1c8d72480d8680b4, 264'h00a866f620640511357b7dd3bc0eddcddcc5a59e9162204c1d85f223ec485cdee2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{311, 1'b1, 512'h21e7350eaa2b2a36fa211d7c6b144fc87b5cffffffff9c3a4d277dd4c34a428a3b35dc4d8c1840740df3876a387e6ae3c97b0a40325ae41007bb1de4338ded6d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00cf3555d277eb8f6fa629e8ed875df1440352e53f32f9509ceecf222c4197c5de, 264'h0084829a1286f98c299ec5c2169a14d0cbf4892a97baca8310279d9b4c98fdef47},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{312, 1'b1, 512'hffde6b2d174d86702f3a46946c7167cabd18feffffffff2df58cb555aad0b0df043b0c01b91bf2ee4827aac1d987f3174e1fce7921c831a0b0aeab1ad1156fed, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00d8dd5094bc40652ddc19d04beeefee8d90fef82628edbc218a9d2de596bb023d, 256'h5c0a46804e7de7c741e5be55a7ebba092dc10a4d1691e6a04ac1690b54acf950},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{313, 1'b1, 512'h55260440dd65e8c48db54c801af143d639f08a95ffffffff9f03419e88a5145c37a3193cc07c160404a9b7d489aa324965d89fc40fab65a71fae34c56afa395b, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h25236b00a0a67e12ea781ae53a929e13c37994ddce784f3c0c33402a43b4a6f0, 256'h117331e5b39fe2a11f5c8bbfa5bb4fdc3659ac0a0efcd03a94362081a4c0e579},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{314, 1'b1, 512'h16438d031fffee5b56365cb1a8f4bc19eb046a111dffffffffc16998d3235c27ddbfe7f1e45105d70ecb963cf511b0e09daa505bc426260466ec6528fd48b88f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0f3564b771337bc8d494a04e4d0518f26d067d07c31689d5e27b503d3652117a, 256'h17144740db21874aa58c0de6a4cadb16c5d9230d4f4607980aabd161d21045ae},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{315, 1'b1, 512'hc0635b12b9164d0a9480ba133839afb60f79f6e7fa22fffffffff18d9363b5c503a5ae2f4cea06d8c5333965149a2cd0ed0491d1f9c8cfbf12fce9914dc22f30, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00bff706d27dc3c8c59951c342244e3c3552216b9225898de130c6a5a8f58eef42, 256'h0e20cb9bffd20d88fe70e5d1f909051528c55efbadbfd7cdcce67de853f64632},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{316, 1'b1, 512'had86d31823a92384efee57d7fc747fc6347312c57d7e61ffffffffbad8263d3a80dcea096adc61333c39ceb1a06bc016fba8beaac8adc0692127ebdaf8bb65df, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ec5c12881dae52168aa635c80dcb0031a43e7d1b76ea97231b819051a861a7ff, 256'h09149c000d1af12d800225c1ba3587a53e5aabd8a8fe78230b1b4c12ba7df008},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{317, 1'b1, 512'h155ee257be62746434e431f20477a5a614b621ca050d7f78ffffffff517e6eeec93db0df6b6358b1f45efcb67e7b201fe4b0f7ef4fe49aed869621bb74d2604a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00caeda2ff27eef0c71a30c277dda128692e4850e589d07f84046342ddaef9842a, 256'h69d422215439150d1da00a0811d2126de5b5c5a85be18fd3c06eb638703e6031},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{318, 1'b1, 512'hde8b1dea4af73e03d31712528653ece2fa048092693f2106acffffffffc4fbe785cc6cb125a5ca069dadd2dd809bc3c6246bc299c2bd84aaaef1085a561dd79a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h3977465917472d3cb67d6fc8888834f26fa47c8d3a2c8e046f70680e3037a37e, 256'h785adced4f3d400b286ad7eb7bdf0b7c0f46d9e7268db5a34e740166caafd14a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{319, 1'b1, 512'h372064a97724ffe3dec873aaa5c4e830fcd9ac84f1c4edb9a372ffffffff621efd798449ba3d7c009467fccb63c6e9a825df2926734122b80e8fc9a6c956351e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h051b252934f1c65f39652a893e9517f049af42259936832cc3f8ff56d7f3cc54, 264'h00867bc57a96eb9d8dc3afd6db11b527f19e4ad8c031134ae6ec9b2b6ee092549b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{320, 1'b1, 512'h0a55bcbb94c925c397b334ec37bd5216789d87fc6589738cdccee4ffffffffbca7bb2e94ddb13839ef8da502b39ac80f25abca143e0add021592ea7a36ce83ff, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0162ba940a75c7a12574736d45d60bbb2c6ce7739b04429cc72352adea4666c3, 256'h4c686aaafb4f3615247ff06b97bd76d49b93f65b5f66c93fc2a8a22246536c24},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{321, 1'b1, 512'hef503ce85b5b48ef35abff5d47345a71aa715f5e8e1568c9721a78ffffffffffe6124c567f2fb5b5f476271da455e079b655dc8c9506b65d9e3c60892984e8ba, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00f74e65ddb41c6c01564b3344fcaa8db2b7b73f8fd156e500865a04826c5e4ab0, 256'h6ec0376675b8c3692f397341269667eadc60696d56d8450ced85a65de9d3cfe1},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{322, 1'b1, 512'h5f3afd4f98713d775d93b166838053fa503faf72cf3c00b3c57e0fe3ffffffff7b74af7667db987c9c205466e00679714af8467254f2e441ccbf1bdb9daad40a, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h0091f3ccfb87b3667bea8c6bb07d554467fbb9a77685a6523da5cf97dfa710e6b2, 256'h5559936f9c94c6e4a97c9febbcb2c1a418fbf9f2933dd64def686b3771dc3fa8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{323, 1'b1, 512'h9e670958749c5bbc0cacb1ee6c38e71eede821d75d84cc2fe1335af9f6ffffffff4e9613cec31f535c4c7bdab269d70a8d4b3bdffa3065d91435a4237cae96da, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h0afdcdcf68669ecc53b019d7adbe8dc943f453b74451335a631a2a3dd5672f83, 256'h77ea833468953e14bd428663eebce4b3cdef41e9821704fb91d1515d20078e92},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{324, 1'b1, 512'h1e77a725c36046bc3bd6ca38747586093510952c0a3390d86b508479c0d6ffffffff25680ce9cd685ebae3cafde6315263f7cf4ea6117ccf870d42189ba3abb8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00a197d8f8fa0cccfa7eccfaea7ca4441bda9789cc3e8d22a1d1b14d6deeb2db21, 264'h0088fb12318d60b66b68fe80834172813989c24901e3adbcd4c73860fa9500bc75},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{325, 1'b1, 512'h59f9626626a34d5491d567d0315894fb702c1d7a2ec677a2b595a772b20d8effffffff20557e965f33f606242a59aea4cd565aecb931664e51fee93a92ccaab6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4b3eeeaf50e9f9bae0bfe64e2776bf2db181ab44c763393136927827f3adb24e, 256'h317abec131eddf2117e27ea2bb4008e8fd0f4a32aa41f74eec7b1659c091fd9c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{326, 1'b1, 512'h001db8dc4aade36062b6ddb62bd342923f537cd35c957b47803909be234a3b58ffffffff0b537f24fbdbfbefce08b061b467fe60e7f86531ed3f54c6e29889dc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h464bdc2db7c5a2745a5d8c96a323eb99c175e0f99baa75dbb9c6d29b98facf3b, 264'h00d9328ca00ce32934b4ed340a6e15236cb16e5364cc91ef5cd6f675e048985bac},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{327, 1'b1, 512'ha05bf269c6959e1000f754963c2ee746346fac0d57bb119d3cecfa3dfe702fef2cffffffffddcffafb72da48023b4eae3593eb7c3c2d758c1c6c5e4dc57d53bc, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h270250c591cb20c7978d9f457104afa7c3484879cfdcf9dc6ac8e785e1fd20a0, 256'h09601dc597c123ed7e76bdbe2d146863bddcf357f9217713dfe1afd8f49891b6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{328, 1'b1, 512'h9695a59c40d735b329f1f9c2ffd974ea8e66af6c65a1f7242e1eb02ea6721f9460ffffffffff9327209276e0633e07c96c9a2950a09411d1eabeda48ba90c8c3, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h729a17311a2fbf9f2325117b2cdac18fd6bbe3db4c5a1bd4e4f4f3d8f3d68dc7, 256'h48dd0269cb216e2792f3b410a781c9b10e59abdc553aae2a00d4038f44a2849e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{329, 1'b1, 512'h521abe64cfe7fa37251542760a99aba478c8b79a5eea4ba1fa859e6dd8bf23196e36ffffffff157c00247c6e0a683044034774f96f67cdea42afc9ebe8d78be0, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h5228f97e5d0dfb62cec6820029175867d7d63b179db3e8a9e7eecd1ec55e0b90, 264'h00dc547d7b7b680b40bcbe0cbf9a2d749787864158af3c0e0f8ef08dfcbbb36f7e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{330, 1'b1, 512'h56f7dac71cfda3cdc27537a7fef1026211918d8041d79637eee4bf44f6fda371a67755ffffffff1dbdc9ce7d24880544364cd8cd5925c287a256383c78631a0c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h21f775d3c7f7fe68e84842b30de9fbe4ffbb4f3324b295591e36e4651c14830d, 264'h00afa24a4cd163042da5f767e7088e6fa03efe039a477fc13f6c23270cda91519f},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{331, 1'b1, 512'hba44f1aa7dbd00300b9d114936943eb2585a2ca6cd8f11fd68794b5adabdcfec1919ade7ffffffff099e11a571237729c09fc81d86398317874c3722999b1875, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00dabec42e9c44f0c230d36c45956cd4a8250f3665b6f291f700e73d06fe203744, 256'h23b687c29e03bc69c5491774588e3c519fa1eafae2ff8ede2ffd4a004e233215},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{332, 1'b1, 512'h125406f9b34e4f63c0a2288bf6166292074a0fed2b2c47822bb885520f2db3e2c58186b926ffffffffee3b259d2c85d9ab10b9f10f7f3cab27a8f528b4a82ad8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h381458d6c40c888bf90aef1428bc968caace553f94287e7adaa48943dc55315d, 256'h1e0e1f75489a451fc7cc4bca61a0a7330a5b4dc4283df68e21798996d8c69bd4},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{333, 1'b1, 512'h46943ed052f77d2e9549dfb8b9a4c779959f7b0a78d6bf2dbde3be53634e232d52a793b7778affffffff162f29721e93b2c9de6629fffbe68596e94b26703923, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00e08881dacd7ad6441f80be1d5510b7e29da4c8504d658634f13e5f3cfcf2a16d, 256'h3792541548f0d891ddf95ee40b815fc3ac160cbfe8cd948e0786db7cc20b38d2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{334, 1'b1, 512'h2b88c2f7b3ffbf92cf6698268ef14cba56c268701a73b30436de1465b85a572363de2fbe10e2beffffffff9b6ad94f832c537e1e40dfd29f836574fecb7dd074, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00a3efb0abc9d76e6601cb23d28b0276293eb8d6f2103d0da7b06a0169db1ea6a4, 264'h00c619ab2ba23b20f90bc815d2fd4c345d0381476b164590cd932b40b2263e4054},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{335, 1'b1, 512'h4e29d13bd24e9f13d5e31ac769469a23d44278a67b110f7bab6095667a3a5180bc8124849e31af47ffffffff94e438c9abcb1301833210026c068417d2da4b20, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h61746df1d5f3d30403f5281767cb6601172b26564e97c35d4c68fb7426db4ffd, 256'h7ca2b0a4fb0d58a119a8df391ad3f2de47cb3b1a8fdf04d6ec235f639fe44080},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{336, 1'b1, 512'h5199a888f66bdde1285c6e1d75e11ca4a6fa67ceafbf32d81894eb60ba36c4786868dcb1384710d5d2ffffffff3d60d7798468aacd9f552c97fa4600343889c9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00ce48fc4bedd4dabacc68f71c4f5b58414e9b054b445c4781cf6d9b40d335b4b6, 256'h1e73b8299579684b80801d2fd70d5c6f9a904ab0735b26d27ff44021002c6107},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{337, 1'b1, 512'h7692bad59be557b4e1db6cf148e5f0ff3c273d29d9017b90c8c26236cf78465b335a40716400ae0aaa34ffffffffd68ebefa85c403e0a25dbfeda3354bcc2a84, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008c936b044cf6dbdbe30cffdeb9eb40b4aa48e697975805dd40455e44fa4d6dfb, 264'h00f03bd82bc73dc7a9d518012f9cab5360d6daa06dd0145765b512263b13c3d851},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{338, 1'b1, 512'hadf9dc5a02f2bf38df234e566f0b5ae3c8b5a20cecc2f8565bb8f756ba59b295004e2ed1807a1e579596ffffffffffac7657366f92a09ca3685510feb2182e3e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4bfaa8c78636efe63915dabaaee914deaaf4a06ae473679160eaeca88d5cc116, 264'h008bc24546613e4811facecf605d6b1f79b442c3d8fe458c1c69334cbee31ef532},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{339, 1'b1, 512'hf9db531c8bd06c7272a9ae2de6b4cac8e0281438eac5689c7f763241db7b88b4a6c71d53a3d03222f6195dffffffff0b690ef5a310f733b13a1bda4fe964a38e, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h130fc664eccece7b71a0a9cadc5369fb5bd54ccc53fd2c515e5ef232acd1b965, 256'h4372a69ef34ec2b296dbe94c5e8a8881645b9c0f6b6c4270c19b81493eb59421},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{340, 1'b1, 512'h273f59b9ed631e0fc10467687508d817c2229d48e45efa2a6783290c6ab048c048a882eef2730e7456b3d4b6ffffffff0369568d9ede46d524123c6cdf78afb6, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h7b675a89f3165e2ad1f3ac4950898d17e7cd869df4ef58aa54901d51193f91f3, 256'h3a7ea099d7c2909ff4a5c3c286d9f7739f38b7e44605ea3f515fde117a4519ec},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{341, 1'b1, 512'he6ded1492cb08b685e2c14f2f11d4bb2fe1601c47019cdd5bb3a42aadbb88f1335fe76ecf455cde30b30e18d35ffffffff921892b8870a2d1248dcd97ed5449f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h393a056a5ce76dc161daf1a6a77afb72cacb809d4173b9126e636a01cf7ccea1, 256'h0859e4195124e11e40db391a7bf04f3ecd7dffe2a5629aac9374468fe8f1701b},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{342, 1'b1, 512'hef9ce8e0e84c667ba940ccb1d3317daddea8b9888a2ef5b718605aeff060c7140522f73cdb7670b0e055a2646509ffffffff81c895857965435d4c4421eaaee8, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2d9738a6e36c24a5dcde61ff7fa5ecb1e96e0077a4a183e8953745cb9461e5fa, 256'h55abb27fad179d132830f7e5dff0d26a63f0141fe2288b9ff7943c3a482ac124},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{343, 1'b1, 512'h388b354799942c6595ba49bc6bf8e7ca5c06c6ae8015c0f58e69192d96cc60e30696c1284ba98c1b22c5c7f23bf8e0ffffffff15f579e355c7258262f0fdfdfb, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h460f528bb6f8adb55626c5166c4572a93c3825dd1a695822a81c9e75e37fe8fd, 256'h0197c8b83193110f0426a417fae7ec3b99fc669371f1e7debbbd3850f6956c14},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{344, 1'b1, 512'hc6bf307fea8c2799ef482911ac86779072e5757f934a3671ad8c5a9e372bb2ec8d318ee3bd0cc4460f9050c937a3409cffffffff81c81c22e9468fd07ec09f55, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2d13939455192c22b1f18f7ca82ad4265ec2c4dbd124ae4a2b0017984512c9e9, 256'h3d9e4fac784be61e2decb75a1f6768af21873eb49881849b936036b19187a734},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{345, 1'b1, 512'hf5f21b002be6b7b3a605b3bcc5a3a12aa0b905565d958028fb8c44d8e5182b6ea4beafe63cbdd96daef63b98ae46ff91bfffffffff3ffcdb29cde67329851fd7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008f2523bbd4a2f4d144c0b7f7b5da84ce20d0d4f551cf5e0ad2b0cb06c6a207f0, 256'h05e46a85f61e1676def59d819220edcdf421db36efbe00bda7f9e331d56e8ce1},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{346, 1'b1, 512'hd88d68932ee321d611334d87de84ef4240025f9d0c8f11bd9aaea2e7729ad87ab0ee66d229b2eb78221050b375a54bd698a2ffffffff0967dbcb983a8f09417c, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4f60878beb2755b35f7152a33e416e16e10f77bca2ad70b09c86eff148ca6fb3, 264'h00bcbc6fa18d8ca570b4a9a5f2a8f6ff9db3e3370ffd3e5a7e19880990f6f8e614},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{347, 1'b1, 512'h611df311628ef69305da2acf952b7289eaabbf389dae756f08c459819db39b7133f02dd126e0442f19bce8ee83cbaabdcd974cffffffffb7195ff14e2d445864, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h009b148c63588ee8f22436a61d52ae8a60c3f35007dde8bb6e31997d99205973b3, 256'h2015548563168f496c7b115bff541fd71fc926448a4554a15f97c58fdd039015},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{348, 1'b1, 512'h4f34828f9520f17da9e588884a26df5ab85e8456184bb19001abc926a180c32a112ba4164e81d69b8fdaaf3c60619a7d1a5840b6ffffffff8748db5ab09c4a64, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h2b7d769ea682af0be42866cf3ad8865b12d4b37c3708fb2ad0dc5c87eda10154, 256'h11d8c48ba6c400f7950f9dfd9ea65617b3765db0e79778bb079fbd7db67b68f8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{349, 1'b1, 512'h4a3d25b54b17b001046f323462e30475caa0fe686e8fa4eaa3b0cbf604de9812e2cb4eafbbe44222356c1e1702c09078e7df08dc98ffffffffff06067e01ce41, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00bfd3ac436e5c4d42f15fbce06d9859ad82d460d322a8c4c1d06ec318fdff4f51, 256'h335bd5d0619a5290c7fce42aaa97ccd52d80528a09a62a4ce8d1e7cf00db7a26},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{350, 1'b1, 512'h6a763ddd1f348cae57162f918abd67d536a03431ed29721e179403366c3fe64f1083d4a64cb7a9fddc7c5a3487675be4078be3b484ffffffff2d5a70dd12c49f, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h56a5c2c2e803e66c5751fe8fb348822609b167478cad4030e7bf6120fd535bb0, 256'h7b3fee66768794c0b362f2d40ad64fdf03e0fb0e8a47f2034167aae2ca383c0e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{351, 1'b1, 512'h0844602883dbcf60972c8b943b5ea020ccb0d19c82eb86cb18d4225a79f97279539214d6e3df6ba6af165c9cd95b8b67a36b39bbd101ffffffff5a9aa9794dd2, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h71bc399e5643a1d8e2afc317e78a2c43d76b6d87f17a5809a7b6d19f922c2e62, 256'h057e7615a2c9033ef0d1a3d3020977002395e196d3b8206c9afecfb98abd52d8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{352, 1'b1, 512'h73672c1037e14e2ed10a0928e8938944667e83879d16f2688f2fe0087494b9f496471dd4e27f5cfddfc4b5efc4e7fcd511d2f67ea879f2ffffffffaebc4501e4, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008f94bcda036e64783935456289aedcb67232932db1ac2e8ad1ca970b14d47a1a, 256'h21a71528f9e8fe6067ca74cc0d8b4b48270aad9ade9db44a98c98182a5e8f208},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{353, 1'b1, 512'h1c28cbb7dcfe2b79763ccf8ebcb7939ea373f7751d8b3965fdcd8b62e8360f619321855d0fe872fcbb3509f48c195d96b1d765983c695686ffffffff51d7cbd7, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h277a0c4f34b2749fd58f55a0f373430f3c868bb1f485d477102b3e797cea5560, 264'h00bccbec7dc1e2740751b7cb8968e7d388e136d7647a29c6845bcf3759f44bf389},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{354, 1'b1, 512'h823e30e3f8bce86e5790d073d931eed5a7ab1f52fdaa4a2522831c73dff05fdcc91829a51c8c0c97c24def713b52643ab17a700ddfa0988740ffffffffca2992, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00934762967efc8c97655cb73d7168d1abb5889e55243dc67c1c5517d6298ce2c3, 256'h44c32fb9d2b5e6f9c38226538776538a55eb1bdfbac44e3e1229337415645db6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{355, 1'b1, 512'hf2104bf641a8b485448e73c4b7de7fc4ec1d3e06eae0f264dbdadb0d514a7aa2ff1567a80e8156c2bd97579eb1467c0efacf0fdd1166e87838a2ffffffffc8e9, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h008f052802126f222ba3ade9cfedf59fc479a120ed8e59366b1be4f3039480004e, 256'h3e14e9209be9dc6d00ed76cddca1c2e5b85f112bffd2779f45f246cb60c319a8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{356, 1'b1, 512'h3db47a2cad8a1c43f31ee677cef231cda0f3853901676c1732771602ccdcc294a38fb8df77d5e6e5737d4c8e05953aeb81edb39a25931717b3c154ffffffff9d, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h4456d6792ff7e4d27517113f309177c26ef3bf6482e131d43f9d8b80e954d61e, 256'h4ffbcc50a7a69dfce92a47410f8574f7b0abfc8b4c7f74ac0dc1c1183d393482},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{357, 1'b1, 512'h6becb022ae22ffc4efd852cec1259abcbd9936403db48920bab66dff9bd34bd1ba5c30d1e8752af80d13d9304dfb864e834181cff7e8be9467cc3617ffffffff, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 264'h00c0e27a8ad306f4ed4dd77edcefb61a6d8f1a9f6546a9969e794432fcb576cd49, 256'h67fdcab3395eebe53dd03b9cadd3eb62d84327de15498b60a60b023fea990436},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{358, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2927b10512bae3eddcfe467828128bad2903269919f7086069c8c4df6c732838, 264'h00c7787964eaac00e5921fb1498a60f4606766b3d9685001558d1a974e7341513e, 256'h504d070e4cf2596e560c1aadc63c573cee0bf8c4d128292c23b47a294c607703, 264'h00f181213b28b921af292ea2fbcb8af4a0e14e2c5aa603c45dab7a46f05bbd5d85},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{359, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0fbf9d131ff8a037747ac23246c5b0e0ce09a905432d3d75477af2d2993b1e0a, 256'h4b14e93d4574fc2a553f85eb3c4c0658a1bd7e1cc7f08d47396e76d6d40ed772, 128'h4319055358e8617b0c46353d039cdaab, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=128b(16B), s=264b(33B)
  '{360, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0fbf9d131ff8a037747ac23246c5b0e0ce09a905432d3d75477af2d2993b1e0a, 256'h4b14e93d4574fc2a553f85eb3c4c0658a1bd7e1cc7f08d47396e76d6d40ed772, 264'h00ffffffff00000001000000000000000000000000fffffffffffffffffffffffc, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{361, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00920945522a364975ffc27bdddd7f01ec26ef8ac48d466a81fbb1d02fc89133e9, 264'h00ce7d01190e815daf1d18e5932ec8a3d83af59c7f66738b6521a9850d794a4ba3, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254f, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc63254e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{362, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00e0ce6d55dae257d10a06be4fb7333e68475407a401de84ff86a931ac022a4513, 264'h00802ca56c9a1d2f67e8a45703b174f0562dfb7e6a532eb1743b3ceb49f9bea420, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00909135bdb6799286170f5ead2de4f6511453fe50914f3df2de54a36383df8dd4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{363, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0c5baefb69764c3a55e9d3ef10a76f652ffa697794ab91169878116d058420e3, 264'h00ccd7b9153694151ee2d05048e40fe072d8e0f481af5d3d0a9e8cf39e1ef7e0bb, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h27b4577ca009376f71303fd5dd227dcef5deb773ad5f5a84360644669ca249a5},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{364, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1a4cb39a674bf0bec4be1a5b035ae18634f4b681a330c1f91b42366a0a7c7532, 256'h0b3f8018da54a8d0db30f7c2b3f04dc011a4a1c383221e52187632a565e5795c, 8'h05, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{365, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1cd72095fd856cf29fafb81c25f7ff24dee34eeaeacc0025d512091b1f1e822b, 256'h427eb3bbb915209e064bfbe1a1798ff6dac8d0add6d753bff4f128fee7e00f89, 8'h05, 8'h03},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{366, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h697cd5856c8c347fdfbca4c2cb2fc1be12f1611f190333b80a5cf4e0f7d48dab, 256'h5d08740936bbc46c90b1da916d5ef39c3d9fb9092f579a43d911472022a7fa90, 8'h05, 8'h05},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{367, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h69d31ff52dbc0935508755cd48cf3f30f0ea78fb670048983be0ebacf4de1076, 256'h773c9dce9aa24b783d8688d63547dc987d4650f20c1179e6ae5d4f14f6d55cc1, 8'h05, 8'h06},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{368, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h69d31ff52dbc0935508755cd48cf3f30f0ea78fb670048983be0ebacf4de1076, 256'h773c9dce9aa24b783d8688d63547dc987d4650f20c1179e6ae5d4f14f6d55cc1, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc632556, 8'h06},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=8b(1B)
  '{369, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h22554b95fcd18cb7cdf7db4a57b259f3d40f5c7cd5cc907a1d0861b3b835fb2f, 256'h63b92993893f14bf17fb9bdefbcbb9404c1985e7a19699d048483702f7e25547, 8'h05, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc75fbd8},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=264b(33B)
  '{370, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2f5c464f48423a87806e88e2e6b4e6f947eea1a5f2c0717897406d97dd3c2865, 256'h61b62e969abf04b840be9587a2a16c0a83ff3bf6812b7257c106a26be2e71d25, 16'h0100, 264'h008f1e3c7862c58b16bb76eddbb76eddbb516af4f63f2d74d76e0d28c9bb75ea88},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=16b(2B), s=264b(33B)
  '{371, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h27527d9ba351f69285cbd9ba144b9e7c6c957d418c8bf63925fb934ab587d385, 256'h216a626307e247c3d5bcf489b52ad4c1987973d7d4cc90fb5b1f488d80134656, 56'h2d9b4d347952d6, 264'h00ef3043e7329581dbb3974497710ab11505ee1c87ff907beebadd195a0ffe6d7a},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=56b(7B), s=264b(33B)
  '{372, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1bfc106d79112f08439a4ffa4e06261bbab3031ff7ed32568172caaeabae2f90, 264'h00b894ecc8922ace776ed6d1526b7771f2cc43b0e84bac400541619e142319059f, 104'h1033e67e37b32b445580bf4eff, 264'h008b748b74000000008b748b748b748b7466e769ad4a16d3dcd87129b8e91d1b4d},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=104b(13B), s=264b(33B)
  '{373, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h71e13191229197eefe9224be11217878635056fd8e558b74121036043cb75017, 256'h09a09bc004ffc98a4051a3fb9798cb9fd5c17919ecab9ff8459a7d561f3058b2, 16'h0100, 264'h00ef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=16b(2B), s=264b(33B)
  '{374, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h15b8867217bf4d531a5618509d9cddc6a3ff4fcc55cc94df82d9952b42ae564d, 256'h7234d5c43238e591501c1fada39a60057fefb46b588d47cbedb529def080fb83, 104'h062522bbd3ecbe7c39e93e7c25, 264'h00ef9f6ba4d97c09d03178fa20b4aaad83be3cf9cb824a879fec3270fc4b81ef5b},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=104b(13B), s=264b(33B)
  '{375, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00e7c1fcc775b8d46770261c413291bc9d913c7785779870eb475f7437da3ee1a0, 256'h16ad8986f7ef63d4237a9c802e5e49471d248e4df64283e77608ee191ec61f3f, 264'h00ffffffff00000000ffffffffffffffffbce6faada7179e84f3b9cac2fc6324d5, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{376, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00cfac11bd4b7aa0a29309767eddd337d302f1f42ccab215171f9622992a671e4a, 256'h1451102ad100a24e6fb5cb130c69de2a61fa50f2d07a099d73ae96f971593588, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{377, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00cfac11bd4b7aa0a29309767eddd337d302f1f42ccab215171f9622992a671e4a, 256'h1451102ad100a24e6fb5cb130c69de2a61fa50f2d07a099d73ae96f971593588, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{378, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00ca99e8cacb96b9b73a7ecf478617269f08971c307aba958692381696c244443b, 256'h5c5df1f740db3016b0ad298997131cea685b2ba405c3b0f722c6992bdaa6fd3a, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{379, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h3c31be015178a9c3d3cae9103bf25bc11a709316d06ab46c01f884a8eb33da2e, 264'h0091f32a1352712508642c4774ea67049175161cb2bafd5524b813274b140f8e99, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{380, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h355d9c3f97a282ac17f7bc98373f271d6a2bc02eb964f13c1e2d7debff4a02fd, 256'h63282e78fb9b88f81413bcf95f16982d9f50e7f94a5d28685b41da997201db5e, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9, 256'h7fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192a9},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{381, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1c959964cabaa5ce966b95acda1c5264847a780426c878d716d73ae6621d3084, 264'h00d3fedfc4f9c3b8cc8bc6539b821ad208ec08d5737aaaf1801d666ddc37e54faf, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{382, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h009842a82a83932d5a44daab14afb79968dd24d9ffc58e638586a90b0f25b521dd, 256'h38b2c05c8d548bcf5ab2a906e2f3fbdde7f0b9bbdecb852297d55ae34257f8f3, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 264'h00cbd25189e59c5c367e7630cbd4c4cb1512c194cadf353d6331f9f57fa81b338e},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{383, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00987a839ec570964d3a1bfc6a0334e7328c1624677c66b8fef3a5e64d1178ddae, 256'h5577dfcd0fe00da9e1d8bb8bbd952aaa5bc10ecb14cae4e3f5e28c506bbc3a21, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{384, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00ab6590ad5134f8e1bf4581cf90ca0398ceb92861c2af06928cc0303d9654ca3e, 256'h1d821f6a357dc173f22a3b77145c057a632bb56f31514e31d6d2ed7fddeade55, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 264'h00aaaaaaaa00000000aaaaaaaaaaaaaaaa7def51c91a0fbf034d26872ca84218e1},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{385, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00cde41230f0cdf732ac76e5f284cb7f46915ed309b48debf245f3ff2f243e9366, 256'h240da36ca5ad289bdfea83213847b14a73079705eab0a2a28aefc999e5ed1504, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bc0f3a265e2136998083451163be66f8b6a673bf5cb08a0e8dbbce4319af6977},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{386, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h36c6faa9f6dca42ea8b0e6d02d36c3941582749251bfa88c35fc8a8e9ad51cda, 264'h00c44ce5f20f36b4ae75cc7291678dbff188cf8c838b8963eeb8b78891795a7364, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h2a06d743967a1330ca91cc46c9394512cc85b4f1b9355eb7f4bbe53a32b76cf4},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{387, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h709e58a12b12034173395bf91e68255d90d8a3a1d5875c75f87787d9a85a0929, 264'h0080e09b79f43489be726a4253ae6c05adce71bcc65389254923cbfacc0775bff6, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h008a457017b290d6edb5455e167b9944f67dc5ba958c7c8108ac56e8596b9bc9a1},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{388, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h0086664a9e09db80dbe3bd0158cc4a64a2cded9c852b455f4443e97cca5569f7cc, 256'h7454f96b52a27a43a1345b5d340902e147880adaf2fe691c168b4203ba2e1df4, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00cbfaf812124638c0b98c18cac3dd8d0848ff921f26aec42a708df7b6a97571c7},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{389, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h623c668c5dbae406e7b4e8e97b2bba2028586f2e3c31f694d9fe87a3de29f843, 256'h3ac7eb04891898dd9077432c38cc978049cab7721630ed033095f850ade83e3e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00af812de3638bfed9c18cac3dd8d087e7350cc7062635266a525bff486363cc91},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{390, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b034897e2a74a787e008b14c62882eaee0e6e53a1c8a58f709a54432713c20fd, 256'h28e07de2ca64b5e215d25d0530d7807df11b98bb39c26a2405388ac0b163fafc, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5f025bc7c717fdb28319587bb1a10fcead32935ea552ae4fb0fe33cdca6473d1},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{391, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h14c4f6210b628edd441651d3cb61a07f7ca87629a9e0add5a4fd92902a20cd25, 256'h5146bebdb22b4d49527ebc90ba6294784ae7ca664724d45a466c9fe8b8699bbf, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00de4130d1ed9120b8c3dd8d087e7630cb9a8402519439af08e96b342788c6e84e},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{392, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b5408eefbdb7480fad4c1735f378c9a1ded28cf476835f27b6fd3b8af5e4c596, 264'h00a60a806e244c63a798baf2fd5a66c6c0d7f77952ba2d74b0fe3652811caac6f0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00ec618e7b1af40be0d052f5a020388fc6cafb822933c1bffab137885f52e89d3e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{393, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00de9e22bc58f4b9c913e7f7c26fcbc5d7f6bdc9fced5f520ac88e8a03290be403, 256'h746a125844509d79840e35440b312dbfdf4ab8ab0011e7c36bc9e01201b1b0e0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00d39813c8102fe0f18cbfac4b0fa028e6e48c093c59ea00dc99fad50f2d614a3d},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{394, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00ee3bfd2e1c3d99acd88dbf6fc9a3a8f5686b50a6a3e9215f57e83a81389836a5, 264'h00f8ebff9a3e463d47ec36259fdde694bdbb880b0a09fe9ac649d691646ba624f6, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00e9fcbcad906698e02d9aba57b3c4e9eefeaf3cec7a980c422fe7f6303fc4a3ab},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{395, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h3c0c4d0ad0848d1335b12a8919d32fafc5f2b0d5c2f3cf6494b06ba8eb17cb29, 264'h00dd7054095454fdb519279cde10259ec5d9e5e4b5a8c4daca649a150f2dbf21ac, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h21f862ec50ef64b3bfbe5d774e20cc838320437725338a3b32fefe3ff159dded},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{396, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6cf91440818ea262b9376e23f7b530b9e44edf5bc6db1a67dd60cc722975d623, 256'h17c19e7d6ebc0cbdc89388242d604ae94ac4ca179ef2cd8bf33fbf738afcb39b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h43f0c5d8a1dec9677f7cbaee9c419907064086ee4a67147665fdfc7fe2b3bbda},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{397, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1b5afcf39888d2da7215f36421a85c4217b0ac883bf5957c2d066efd8bc89f18, 264'h00d8fb3b6aca0b3577a883948e016905065a3fdc13d6f433172ee0f16784e52c78, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h65e928c4f2ce2e1b3f3b1865ea62658a8960ca656f9a9eb198fcfabfd40d99c7},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{398, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00890d36db646c27c2e6c7bc7fdc3f0cbf66fab36d13279b9ecf6e98457d8cf492, 256'h07a83cfda8e9d0375404c6cbff66792eef97220239254000b4bf983e6bae26d7, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00c522b80b59486b775aa2af0b3dcca27b1d565aa199ca0fc6d008598e33ff7779},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{399, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2a1571ed0ffe39574d030b406f638bf88eea5b4b50754e93431fe0172fdf2fbc, 264'h00bc77f601dc6dbc88cc2b560e8cca5e738f2c769810b2c8762dab917adfe24535, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffffaaaaaaaaffffffffffffffffe9a2538f37b28a2c513dee40fecbb71a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{400, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h612b4467c8b3b8ecbf5374997ec7db8cab2bda9e431982c49727f3fcefb10b47, 264'h00b9d1ecc026c3665425730128138c4e181c61ec28b38910ca59e5fc496ec31f08, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00b62f26b5f2a2b26f6de86d42ad8a13da3ab3cccd0459b201de009e526adf21f2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{401, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h34191b6ce8865c2230a514b61e2b2730c94beb072e9de309872aea3743bb3e27, 256'h22d202fc59984e7421a25e6a82664b5080f72ab28df9c0af4e1e300af11ae9b0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bb1d9ac949dd748cd02bbbe749bd351cd57b38bb61403d700686aa7b4c90851e},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{402, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00d533c620a8fd3d5a8342caba89eadc25907d1e9b6fea48ee8f806aa772f0c80f, 256'h70e09c022fa1139da32a456ec024949824477bf0bdbf603e8faccd6b205d263c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h66755a00638cdaec1c732513ca0234ece52545dac11f816e818f725b4f60aaf2},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{403, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h0091014bea8705a022972e12b176c96e84c0b61c05eb1c6f8c5c1db731d54d67e2, 264'h009060ef6c764d8d47ed5ebf8f6c23835cb89f8b056cdf7e457f9273b6477ece33, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h55a00c9fcdaebb6032513ca0234ecfffe98ebe492fdf02e48ca48e982beb3669},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{404, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h287a7f8edfbb55cbb56d6b7be5b96c410a85a35bc6639661a92bd653e1f59688, 264'h00bbd133a77828493b3e0f867f34acfcac099415399a6b1106a0f9420c06f8bf94, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00ab40193f9b5d76c064a27940469d9fffd31d7c925fbe05c919491d3057d66cd2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{405, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h0082eca524c9ee8475ec8948721a9409b5090c6c28866d0c12669bd5cb7e685a58, 256'h066b1e7135946a425ddd228076ea24d131b9bd2eae6b51c8083857628f260b80, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00ca0234ebb5fdcb13ca0234ecffffffffcb0dadbbc7f549f8a26b4408d0dc8600},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{406, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h009cc512b58d5b921f91075441b0df61e0381459de703a84523cda31dc18549ff8, 256'h5647dd4bd39f6761a144d81ef39db7bc0dedbcb15bdaf084e3a10fdd10bd906a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bfffffff3ea3677e082b9310572620ae19933a9e65b285598711c77298815ad3},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{407, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00aa9d33c76ccd011ba23047a420840374b4fa3be480c65263d543baf2ccc6141e, 256'h5ed3b42ad9527869fae92914b82b952d2c31c8fcc85b4c100983096694285766, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h266666663bbbbbbbe6666666666666665b37902e023fab7c8f055d86e5cc41f4},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{408, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h2812996934db1357048a1aacb07cb2a8730fbe530984a7a5166f84748ff63e4c, 264'h00e6e8a80e235e216e1a9e75ba3b3a321af51d2e4524ad3c8be99288463b91155a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bfffffff36db6db7a492492492492492146c573f4c6dfc8d08a443e258970b09},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{409, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h008286d34afa1904ae756d73bf02a6b6a9db1eaa1b8351ad713a786dcfb829135b, 264'h00f97922dfe80cd4f0e438a8d842e7666853436d972860f715e622a1e876db4251, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 264'h00bfffffff2aaaaaab7fffffffffffffffc815d0e60b3e596ecb1ad3a27cfd49c4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{410, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h4b7b9990a6c2c5a810107c09ee09cf3388c1a6e82aaa44c378d9886e2508c2e0, 264'h00867e7632fcc312fcfdc01fb6a579ce6aa6285563b1adbb3272f0e122f9de73e3, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h7fffffff55555555ffffffffffffffffd344a71e6f651458a27bdc81fd976e37},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{411, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h568426540e19be6404e6cb4745fc7a943c0c059d7c7baf3bc4fc782e9aedf2de, 264'h00ba7fb20ad12a886c53945d3cdb019afa8b0d58ed307d55f556acf79ec89012d5, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h3fffffff800000007fffffffffffffffde737d56d38bcf4279dce5617e3192aa},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{412, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h1bebc1a6823107d1263219e36d2ec1957d20b0b450b481c9de46ea9294d48b66, 256'h72b7a811af9528e61199f4a2a7f30d8685f5a04767b59276e65a732e8f3950a1, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 256'h5d8ecd64a4eeba466815ddf3a4de9a8e6abd9c5db0a01eb80343553da648428f},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{413, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h08a2b7fa625f09106a1a8d98f831e53d918fb330d6c388a7b80df98bb9e9c934, 256'h478da818b4d94082517fa9635a8aa5be05323de604fcfa97bc3a1a57a5e80c34, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 264'h00ae36701f241f6073608b5f77d9039a9aec44aa5a12a99227fd2911b001915de2},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{414, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h08a2b7fa625f09106a1a8d98f831e53d918fb330d6c388a7b80df98bb9e9c934, 264'h00b87257e64b26bf7eae80569ca5755a41facdc21afb03056843c5e5a85a17f3cb, 256'h6f2347cab7dd76858fe0555ac3bc99048c4aacafdfb6bcbe05ea6c42c4934569, 264'h00ae36701f241f6073608b5f77d9039a9aec44aa5a12a99227fd2911b001915de2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{415, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h69aac6897b0457e54cac25f24590be255d352a20055004e7caa7cbb430b3c90f, 264'h009113bffe220db9143e38514da0481df67f1717c58aab1a189fb9d4f6e53c3900, 8'h01, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=8b(1B), s=256b(32B)
  '{416, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h449ff6ddbec4bf9bcc3149b8dfe480f9a677c3b8e203d272f3e0a2cf90a2cea7, 264'h0087fcbc0799a9323da3f7fddb4818b89b1d97b32b962e1b3edad2fbed47b58d41, 264'h010000000000000000000000000000000000000000000000000000000000000000, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{417, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b282b1b5bc00c2bb18f28ce678e1cd48c8ced8335af5d8e4abd3d7a7d3616f56, 256'h3d47a55ddc11e966fde2bd87b028e62fc8133def824e3e00528f2442908fe84c, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aa9},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{418, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00facbd6f5e996284a53cb1ca41ffc4eb0a3fd73b73c730194011169b9ada14519, 264'h00c5491ede60614d823b491198df7bc6c6768e064e0e43b7f053ab8f279cd4f4ec, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{419, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00a011801d52a75f4841e40240da49dda8f38e868b4e6f941f77ca9b86665ad5a7, 256'h4751eabf00fc2a7a863fec366975edbcd4885693022cd755c0d8936e660d61db, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 264'h00b6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{420, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00fdfa5d35e42ef91b1842c9f28aeb6c68bd7732935f748168deb718e66608b980, 264'h00d6f85fa678df3cabb55b5002e63b55d7cae11e89f74940b7990a3b167dfa191b, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 264'h00cccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{421, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h0754de71bd21f14f4927bdab77efc57f148b36275c305a86c1d7a0dcfd53bab4, 264'h00989fc99bc725da84197c2f284ecc6030489eda77ef92f8680130622b631af2b3, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{422, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h008aad84fd5d52afd531f1068fb7a10bb365faefa89975597187470d04a8c9c8b3, 256'h27258e32d19cd58ddfd35bd7ea1f063c77c61b7879451bdd3e8f44cbf40241a2, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{423, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b4a01ec7b10acff3dace05222fae05c75368a375d8ce1faf4a1b2def1ab715ab, 256'h61a6642e82ff950f373ace5c0cc298639ab9ae739e4614a93fb1122ee16d922f, 256'h7cf27b188d034f7e8a52380304b51ac3c08969e277f21b35a60b48fc47669978, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{424, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h4efc2bef42b11e0929edca3b025f01b1fa37aceef4cd3e8c2d4beab500856af8, 256'h7716828fc1788c881ae39f534c3e270ca869a578210b5dad8a8938691d0c4b73, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h555555550000000055555555555555553ef7a8e48d07df81a693439654210c70},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{425, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h4606b9fceecc47babcc78de73ca55672f09930aacd560db0a2967a99ef8a595e, 256'h612a050025785c0e7c7763db0bb53c48b6ff0ed1dfb6055df90299e295092990, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b6db6db6249249254924924924924924625bd7a09bec4ca81bcdd9f8fd6b63cc},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{426, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00b6de6de267720d16bccf71fdbe07ebe5c1149f8cfb2041b1d6cabbc9b6656d68, 256'h2d3e21f4025ddcacab035b5da6310361102079f1b40c1ef7c7b88427694c11c6, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00cccccccc00000000cccccccccccccccc971f2ef152794b9d8fc7d568c9e8eaa7},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{427, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00efd3bd1299d4b2bb0afbce2afd90792d8c72e1d29c6092e4681540420664e275, 256'h390a4dbb20d10f7360c5b794564dcd443bb1df94bf6b1f4be5909a22a6a534ba, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h3333333300000000333333333333333325c7cbbc549e52e763f1f55a327a3aaa},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{428, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h00dae9cf165867da6482ede84bfc5b94375529bcb953f26d0cd68fc877088f78d9, 256'h51cadc9f61c55f8e2a04dbaae1251fd15cb12df9bcd072a51971127eaa6ce612, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h49249248db6db6dbb6db6db6db6db6db5a8b230d0b2b51dcd7ebf0c9fef7c185},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{429, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 264'h008418924e94161d350c9fe8dc1cc087de4b4491d0bc694a6862df4e8a555f9afb, 264'h00b0b391af97b0dacbdceb7a982781d0090978efbf76b8e6914250e92ade9a6126, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h16a4502e2781e11ac82cbc9d1edd8c981584d13e18411e2f6e0478c34416e3bb},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{430, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{431, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 256'h4fe342e2fe1a7f9b8ee7eb4a7c0f9e162bce33576b315ececbb6406837bf51f5, 264'h00cbd25189e59c5c367e7630cbd4c4cb1512c194cadf353d6331f9f57fa81b338e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{432, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 256'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{433, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h6b17d1f2e12c4247f8bce6e563a440f277037d812deb33a0f4a13945d898c296, 264'h00b01cbd1c01e58065711814b583f061e9d431cca994cea1313449bf97c840ae0a, 264'h00cbd25189e59c5c367e7630cbd4c4cb1512c194cadf353d6331f9f57fa81b338e, 256'h249249246db6db6ddb6db6db6db6db6dad4591868595a8ee6bf5f864ff7be0c2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{434, 1'b1, 512'ha69f73cca23a9ac5c8b567dc185a756e97c982164fe25859e0d1dcc1475c80a615b2123af1f5f94c11e3e9402c3ac558f500199d95b6d3e301758586281dcd26, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 264'h00ddb577670d5a9b93666df2af7f9baadd8256fca0c81deb2d5cd7301a4b39105f, 264'h00a2bcd9f6228a0aa0a4f066aa674b9b08da252b02a77fd1b2f7a2d85929e8b491},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{435, 1'b1, 512'h86fe1b4ea7ac8e339d04e40087534c61e245dd4a0c22754a0622642bba56de900b2d431e859a36b1a5ff71aee560522eb0d3251e018c2cb6a10b82031cfd37f2, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h532d672c307da2891720d11422035ea25771f4fce0dc9948d754ca4f66ef36bb, 256'h4f296181799d3e6780086d6908ab8642711bd406e481b0ce3af1c44b9f098496},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{436, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h1c58cde69ddb363e7a6d2612771b3e713be8bed07f37bcda4875f152db2ac1ad, 264'h00a66755b078262b6b0d90c74aee64522104aa58b5f82fc5ba98bcef5bdb9d43a8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{437, 1'b1, 512'h7d795fe6a97761d89b35f64e09555951f6ec2a669a9fa03481c100ae158f183e2171e142437d2c3a42352108a22a7e3d797beaf6c3075db419b6f4acca479c83, 256'h04aaec73635726f213fb8a9e64da3b8632e41495a944d0045b522eba7240fad5, 264'h0087d9315798aaa3a5ba01775787ced05eaaf7b4e09fc81d6d1aa546e8365d525d, 256'h6637f14369d1dd112c5691969fcc867e64bafb1f5d8f917a9acf8ecf1dc95754, 256'h457b4a8bdd1c047b12826897991241700dad09666b4f410a56993023b098fd1e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{438, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 264'h00ef9a4672e0a07a0efd5936a77f4ea0fcd69dae6fd95ccba8dcb685e7490623c3, 264'h00cf135d42f5e379f6ef94b6a493db01c740f441ff5b2475638b6b081f445b17e2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{439, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 264'h00b8cb05b278c15df7c6a311b0ce7bb5598fe3a95fdb57683ac0821aa2f5d6fa18, 264'h00a9dfa1cc0c9ae0015ae2485f22ed6b0925e82d96ff695b8c2ed593f02719f30e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{440, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h4f337ccfd67726a805e4f1600ae2849df3807eca117380239fbd816900000000, 264'h00ed9dea124cc8c396416411e988c30f427eb504af43a3146cd5df7ea60666d685, 256'h2fe6f2aaed0eb760223e8c580363630d3041614806e7fbc863405aa4d98825ee, 264'h00f5d2c396e45d9af9fe1b06b27f0db4d9ee66e1855f4846dae5db6b3d8afbc4f8},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{441, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 264'h00fb9e312ced9f95c91248bae25056b7bbd84a05fc92acbd304269a1269bbf4f4c, 264'h00f31426a809ceebb369278a5182bce94835f066cab8654f8bd2339595844244db},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{442, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 256'h284fe5f1c86a55fcb3c27a12d82d794eab9a0d76d1fdc4f25df5a9bf52e8e768, 256'h7aaa75e5a7948be66f06ce52fc3e4916fc93514b08c51f84b73839d2c05acf58},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{443, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 264'h0084fa174d791c72bf2ce3880a8960dd2a7c7a1338a82f85a9e59cdbde80000000, 264'h00812950449ab90351ab0f124774a2633625d0871d42a69d2e473d8ac118b506a6, 256'h50c98878c3699c34f3049e6f9496e3199fb5d860232995205f1761c000af4e07},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{444, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 264'h00eaa4f3a8805c60cff74cec78c6b7cea71ef116c333612a6e0096a4c42450936b, 264'h00fbb3508d6692b8e0854c1a1749ea065262bae7c8b831ece895a1eeda01cebe7d},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{445, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 256'h3d0caca44c21d34cfdcfb00098c95203e08847f4aabab5ae6ea7f365aefbbcf8, 264'h00bb99be729e51cfd167dad22182383314c9d85432309cbe36f4b1eb73e776b249},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{446, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h3cf03d614d8939cfd499a07873fac281618f06b8ff87e8015c3f497265004935, 256'h7b05e8b186e38d41d31c77f5769f22d58385ecc857d07a561a6324217fffffff, 264'h00e4f8b27c3c2c5cb2a6cb9c2049011dd1060085c6e2a15380bcf5224063d3ae08, 256'h4b3a19f1be945cd649f34d965e7eecac0a05ac8030b7cd2d6bed84086fda567e},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{447, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 256'h670ce60d0fc7224c8d06f3b01c4416ee0b3ac12f0cff3e1ad214898389ebc819, 256'h45da7b6fc8f4f766f82c5132735f2ed94130780b444e2e10c1484d5e45f64332},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{448, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 264'h00a22928b3022fd554670a86ed519a48d8448dc90856e9c40589076baff591e076, 264'h00b4005a89aef027e5063a89709fbc66a05eb12d8d34af84f35ea7ac93f7bbd40e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{449, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 256'h2829c31faa2e400e344ed94bca3fcd0545956ebcfe8ad0f6dfa5ff8effffffff, 264'h00a01aafaf000e52585855afa7676ade284113099052df57e7eb3bd37ebeb9222e, 264'h00a277181e641edafbdb359801605791c833ff3b462dac3c4d3608d479c98090ff, 264'h008b2ad68880cede2290a996fe5b7003610c5c9f53e1dcf2cdb2ad815e2ba5c1cf},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{450, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h760c487841a7214e9850b5569d99fe3ff9dddc41dee7313a780921d8d3657b16, 264'h00b99d63e3cc81458801d5fd5926405d33b894e0f96a85c3c4a929a45c828d76d0},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{451, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 264'h009b7e72ac454505017c5377b2c379f31a7a0268b739fca4c97dfe1c9aa4bc548e, 256'h1e65cbee69a42ab0a7ae50e9acceaa0971574fb604958876ad6316c39eebdd96},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{452, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00fffffff948081e6a0458dd8f9e738f2665ff9059ad6aac0708318c4ca9a7a4f5, 256'h5a8abcba2dda8474311ee54149b973cae0c0fb89557ad0bf78e6529a1663bd73, 256'h4a7e44e4a8a9fee22647923eaee0368b3fa408edaa19b406507309b13e073855, 264'h00fd8597585fa0270c8cdf855a7a69a843eb28124ecf90ac53a58a847c7b43c7a6},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{453, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h4589f0c24d1b2f89c2e806f667297c844c63330d6b9a079b2bdd2d95247e3eae, 256'h75daa1da09a3f1ed8de1aacc7039a721c46f9ebcd4672750f2fd9c2f70f1e6ed},  // lens: hash=512b(64B), x=232b(29B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{454, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h377578a81da586eae269f05c9bb2280a517ab3184e02179aca5d64dee1a930c7, 264'h00cc1735efd4b43e8bdba8c1b44f9ec3e62577e5f4f6543051467bacd9eaaa4d4a},  // lens: hash=512b(64B), x=232b(29B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{455, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h03fa15f963949d5f03a6f5c7f86f9e0015eeb23aebbff1173937ba748e, 256'h1099872070e8e87c555fa13659cca5d7fadcfcb0023ea889548ca48af2ba7e71, 256'h7f722716c279f3d14563fbd8cbf3abcd51c3305795609e04c8ed7ede12ae2518, 264'h008a996a370679c3ce6232244d64481e96e47bf6611aa5490000c0b1dffc231aa1},  // lens: hash=512b(64B), x=232b(29B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{456, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h2f11d967790dd4387a218929b3fc0f130238ec6fd9321348fe631a1e607bd742, 256'h3b52a42606d0daa135092d89ab74b3c4e72b4ed213137406d4b50fa84c4ea049},  // lens: hash=512b(64B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{457, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 256'h192d299e96272a0c49ed1b15f9047b54b4878eaf350a7b2f5439b1e3c83f9703, 256'h26513e9cbbaca7946f3d6d90b5cc65a985cdfe089734f944ab74842a4dc4127d},  // lens: hash=512b(64B), x=264b(33B), y=224b(28B), r=256b(32B), s=256b(32B)
  '{458, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 224'h1352bb4a0fa2ea4cceb9ab63dd684ade5a1127bcf300a698a7193bc2, 264'h00ebd7a6f1450f8bb9e9abf9f66c4143d28c8c845b2e260ab0fff3f7ba5837f944, 264'h009928afe57df6b8c90b7af7c3da981b71db6ae3a5a21a4c5a48b71628e5811a9e},  // lens: hash=512b(64B), x=264b(33B), y=224b(28B), r=264b(33B), s=264b(33B)
  '{459, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h37fd00b14ff469a8bb4d2f9c6ca228c4c24b85719389a46099653c41174e9afd, 256'h5f64dc68893cf3186df3e83af70e96e9f2103d25b8ddffecda96e8e9181619cf},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{460, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h3ce339a63ea4cc1a6b12d1e66b91205e8af530eebe3208359c5327b242b2b669, 264'h00f2b1d6dae62bfe9c44b1cbd56cf0de865a1201c0486d658da5fc029ad47b917e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{461, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 264'h00bcbb2914c79f045eaa6ecbbc612816b3be5d2d6796707d8125e9f851c18af015, 264'h00fffffffeecad44b6f05d15b33146549c2297b522a5eed8430cff596758e6c43d, 256'h7bf225bec33ce7fb4014097e350c1504d3374028cda8f6fbbac4e0fa5319a048, 264'h00aaa45d54eba6bb3ce00ce8e63de24dc7ee19069062e8d340663adcac07f097cd}  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
};
`endif
