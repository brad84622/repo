`ifndef WYCHERPROOF_SECP192R1_SHA256_SV
`define WYCHERPROOF_SECP192R1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp192r1_sha256;

localparam int TEST_VECTORS_SECP192R1_SHA256_NUM = 62;

ecdsa_vector_secp192r1_sha256 test_vectors_secp192r1_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'h508423e042b52945e2198ae8b4a97d3810961d886c6ce1e4},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'haf7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{118, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 0},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=0b(0B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac29486546},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=8b(1B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'haf7bdc1fbd4ad6ba1de675174b5682c7ef69e27793931e1c},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'h508423e042b52945e2198ae91aca8501fc2a53d6b79ab9b3},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{159, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{169, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{241, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h1c1af41c461fd2e7ac90cf03775430863e0625609392d689, 192'h56621316c3fb0fc17d1e140c87a8d25141ead133b66fb543},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{244, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h1eba3835f014e1c0173cd60a053fadc9fc0e7709919496a1, 192'h64c7d823cd73423b2c7966c0b248a65e53aaf80af0ab2b50},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{254, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h125b39558823f19874183fc6193c50e4f5fd7f87561f43b3, 192'h1b164d656157ee6fd5c6ed20276f2f9e8e78f40056f4c917},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{258, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h4d23bfb770d8b60bb7ab1aa45e1f6b1da414945fd52215bb, 192'h2d2c57ee3fc517793470f61f38e1ac5dc9cd88618d7f2782},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{260, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h424d505066afc412387b147f0cf96e1ebae3a16f0c0d69ef, 192'h446975a09f8d9c20d2704196f1446f354e79ff3d308c7e48},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{264, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h31cdf0bf4b77c10f5f11bb2ab2a3c778059e076824146523, 192'h058c3be3e7d01be17f1d135745d581ccfcf03ae0ab6226f9},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{267, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h0a666bbd50d32922eceb07fd63971d6b44c06e39f6ae37ce, 192'h13df79819941a6413a4f3ef6f1b62882ecc88b30b041e3ea},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{268, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h654c558777a4fa29fc22026156220258986a262ac65dd8ee, 192'h608e8dc90e569b3d182a663e93f740ebc9fc7b9cd5112879},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{269, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h3247b2b9f8f59df93efea88267609d8a8f7c45a216a2ee20, 192'h4212ee42824f30fafce4fe8286b69cbac02192fcee13e32d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{270, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h37479876e1e96c7ad149ec7725e07ec16ce30f4a849d2471, 192'h1dc2e3642b717b8d1b73b9cf94d8ff070c0b7eed4141f0ff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{273, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h5968579514668883386e05d6d5813f8e3ad54ab595fb51a6, 192'h35006e924c80a145666bb097b9ccf6bfa1650d7b005869e8},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{276, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h193f5680cb656c321307f0cf016c3647d9daba2fdf847f79, 192'h167304e7d677d139103edbf6d09a4291aecb6e05719158b9},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{288, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h634dbc50a74338fe4d0e187111eb776f88a2b7034b879dab, 192'h4201e22c4a85b3232f21ed346ac335e069b610163fdff242},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{291, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h314da19b75e5f8116ab7c6a671e7dadb379a8e86c7452c7d, 192'h6cd48d19c8667db383385742ede00007e484825f214065aa},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c422742cb5d7f990dc9579e85a0339da7ecabda11d7d18eb, 200'h00f547da5ec37681ce86916fc7ef4e91b76aa2073f17531cc9, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h73e5f9eaf96c8c84c93bd31bf65daf4ed20ea0ef67ae0bd2},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e70f06da0e6036bb0ee47fe47836a0f4382e3349ff927112, 192'h6feeb50ab0f618a5557e488bace8fa2932fb03009ed622a0, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h41a92de5298636d693e86db59b3ed26215e70ecfe43620d9},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0094e936a4149ababae26300ec4c915409f6bbcbbce94611d3, 192'h5f326034990f7993559d97901e7ed1808587378cdb236c07, 8'h02, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00bb41507556b67368feb9978e7879305e4fa81beb2c95ad95, 192'h5d7f0e5c3966ad5fee2b5901cc3dec4190175246935ca993, 8'h02, 8'h02},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7e18073ab95a26038e5f35a805c76c8b880f9d175793005e, 200'h008be399eddfdce76e1a42ba16d065bc7186c08b32fcafdfea, 8'h02, 8'h03},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ebb8328e0c8bac41eaf502dfb9e5f5d57014c7ea842b6617, 200'h00c7b6fb10434359da7a29ae458bf2b03b7c9290f79c4196fc, 192'h555555555555555555555555334a52bcb179433b3c460d68, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=8b(1B)
  '{311, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ebb8328e0c8bac41eaf502dfb9e5f5d57014c7ea842b6617, 200'h00c7b6fb10434359da7a29ae458bf2b03b7c9290f79c4196fc, 192'h555555555555555555555555334a52bcb179433b3c460d68, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h73761b8c8aa66d47c302a1af56ce6e64c139de565a2de1ec, 200'h00a526726d7552e162df2c42a7e1523083e150be83167c334f, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691418, 192'h555555555555555555555555334a52bcb179433b3c460d65},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{313, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d7bc9b50e8bff4bb2c6c8116a25a973e95717fd857fad573, 192'h3eb089b00237660aa485016da2f6c3bdec88cc1cdb28eb56, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691419, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691418},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d02ae497238e2def130607b98eed7693a2f8ad4f9294e3cd, 192'h5d8fed9551ff73ffe0d3877cd364ffb104690052cbd0f7e2, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691419, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691419},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4f9a2b948e4ea950a2ec9dfda5ad1b9b619f9eb678b27cd1, 200'h00aff08eaa1b956963e6af3d61f2c5812ce50145fdfe74c2a3, 192'h555555555555555555555555334a52bcb179433b3c460d64, 192'h44a5ad0bd0636d9e12bc9e0a05bc56531434e1ee89ab1ba9},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4dc27b674729ea276d1f9c9b031f2db841497db7ce50845f, 192'h71838b5b21bfb0b238ea9e209ff89c88f8d070933d7f5531, 192'h555555555555555555555555334a52bcb179433b3c460d64, 192'h555555555555555555555555334a52bcb179433b3c460d64},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5a6289c4fb18c344a4edcfd89105c62ffa20cba6814e74b9, 200'h00fd11db2d30eb3b9edaaaead049e57868be475208052a0da6, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h68e686f0eccb840bb80bf08e2ee70d64264fd5162fe2159c},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e8955850e22d5c08c319b66b9abf74387fe6d209356b671e, 192'h3cf26e4a6a6df3ccf2aeb15a3d949d382a7ef87cbbc419ca, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h7d583e05abb0744a5ad0bd0604d88c454169c54db223a428},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ac3b619c03c378e6018281e70138fb656d9e79c14287c223, 200'h00d7368c53015b87e03dd88499556ab89406e5928f90094395, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h4f1696d5ba25729655f53877ae5a3c4631776eb4bad5d13f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00caf74fab27fbaf4c4a1da037583d7c3ac651df9863d4c4fb, 192'h21d54ffcdb5c2cc0790c712de4d889febcdb49fe890315d3, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h16e1e459457679df5b9434ae01e9721bb166f5fa2de3b3e3},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h3f0635d2d1dc63d37a911bb0b5c4afea9fe2a6f8243ab27d, 192'h6178cda8f95d86e2f8927ce903ebad88e944a07ed8ab3417, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h347343787665c205dc05f847177386b21327ea8b17f10ace},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c36e6fa900dacbbcb6aaca3aa6efc49b453b1bd4b04ce158, 192'h2e351f235b2f2f66a9383597c10fb311572f011f52bc0902, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h3561529936d8c7ffffffffffeab455eb8a9a41f7f1676529},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{337, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h2de010ef4508cd806b145061f5be2986c12fd98431f403ea, 192'h71037bc5d2d3d3e686518cfc719bd2c00b19027e7f3880f5, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h6ac2a5326db18fffffffffffd568abd7153483efe2ceca52},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0080ed329fcdf36f7f8a33ca2bb65a71f52864d75435b0e7cf, 192'h790c28f5a4e82c9ed3a3845799ee4dc6426cca1322db7d3c, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h29936d8c7fffffffffffffffef69e514dfd0b9ad6b3f3dfb},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009e74033763a653ee1eb69584268de7012905f003869a52ae, 200'h00f47afc4fb2fa6a3f1572f165ffe998e40ed5125b83f51a5c, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h155555555555555555555555444fd40903674c4848cdb15e},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{342, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h31d49b617bbd70c6177bbdf7bd7d48c4b04d3033ee2428c8, 200'h00f9032538ef821c03f6cb6891742eebfad72d45fce55fd5e8, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h2aaaaaaaaaaaaaaaaaaaaaaa889fa81206ce9890919b62bc},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{343, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c1f93e227ce3ee8dd56a70e8825b2494c244e1c7c5876e10, 192'h185684cbaf96e3a47302319971ddb1cf52073dc0a2324565, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h3fffffffffffffffffffffffccef7c1b0a35e4d8da69141a},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{347, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0098764a1282d3a1efd6e412e205a226a52c91200ff6728f76, 192'h712f8b75ef23d945288be4b6af16d1e22fd42bb8a8ff64a6, 8'h01, 192'h555555555555555555555555334a52bcb179433b3c460d65},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=8b(1B), s=192b(24B)
  '{349, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009826be07a2fb115616e96e29a35f663c45aa6aa44acc0d2d, 200'h00ba68408829c30e55b035719117565d40e3ea8ddd656faa01, 192'h555555555555555555555555334a52bcb179433b3c460d65, 192'h3333333333333333333333331ec631a46a7bf5238a906e70},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00eced81c0c456fc3238d08f92238962778b85bb596b27768a, 192'h14b06921bb4656b7e800d4cf98d06f5b381b8aa0d7fa7ad4, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h555555555555555555555555334a52bcb179433b3c460d65},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h37697388bfe2dafa44b03111fd3f9de97664e109edd25f76, 192'h59445a4f6e038cf3f541250ca40a89ce7d3692c9fc0e0975, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h3333333333333333333333331ec631a46a7bf5238a906e70},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00dfa930300cdc9ee289effdcc06c26f332b6a0ef598428495, 192'h4c2e5626703904f5643dc693062c71995e789f9c9663e8b6, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h6db6db6db6db6db6db6db6db41f1d8172d52c42796a335cc},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{361, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7bff39306ffc5cc10f34609435ec21eab7a3b49967f7f3b3, 192'h6c0b9346b2c981d59f77079c8f53923c496c73f7ad7d07b1, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h0eb10e5af0643b62b86dc5451543e9035e00a5276c1f7a3e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{363, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h07192b95ffc8da78631011ed6b24cdd573f977a11e794811, 192'h44a5ad0bd0636d9e12bc9e0a05bc56531434e1ee89ab1ba9, 192'h24924924924924924924924915fb4807b9c64162878bbc99},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{365, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 200'h00f8e6d46a003725879cefee1294db32298c06885ee186b7ee, 192'h44a5ad0bd0636d9e12bc9e0a05bc56531434e1ee89ab1ba9, 192'h24924924924924924924924915fb4807b9c64162878bbc99},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{367, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 192'h2a551b5a39771e436de636d6259ba6afb1afa5d4d897ccf8, 200'h00bca9a6ea5d92d656c4ba4f2dd85c9d86d0e2445fd5db8692, 192'h1c5298437de413483c777e1133e62d5b81848747b89480bb, 192'h03b56152e323216bd9d9e403c8cd229a68014f6e2b69015d}  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
};
`endif // WYCHERPROOF_SECP192R1_SHA256_SV
