`ifndef WYCHERPROOF_SECP256K1_SHA256_V1_SV
`define WYCHERPROOF_SECP256K1_SHA256_V1_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp256k1_sha256_v1;

localparam int TEST_VECTORS_SECP256K1_SHA256_V1_NUM = 132;

ecdsa_vector_secp256k1_sha256_v1 test_vectors_secp256k1_sha256_v1 [] = '{
  '{99, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h00813ef79ccefa9a56f7ba805f0e478584fe5f0dd5f567bc09b5123ccbc98323, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{100, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h813ef79ccefa9a56f7ba805f0e478584fe5f0dd5f567bc09b5123ccbc9832365, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{104, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=256b(32B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h813ef79ccefa9a56f7ba805f0e47858643b030ef461f1bcdf53fde3ef94ce224, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7ec10863310565a908457fa0f1b87a79bc4fcf10b9e0e4320ac021c106b31ddc, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{159, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h900e75ad233fcc908509dbff5922647ef8cd450e008a7fff2909ec5aa914ce46, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{180, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{182, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'hff},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{293, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h28f94a894e92024699e345fe66971e3edcd050023386135ab3939d550898fb25, 256'h32963e5bd41fa5911ed8f37deb86dae0a762bb6121c894615083c5d95ea01db3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{296, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h325332021261f1bd18f2712aa1e2252da23796da8a4b1ff6ea18cafec7e171f2, 256'h40b4f5e287ee61fc3c804186982360891eaa35c75f05a43ecd48b35d984a6648},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{298, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2bdea41cda63a2d14bf47353bd20880a690901de7cd6e3cc6d8ed5ba0cdb1091, 256'h3cea66bccfc9f9bf8c7ca4e1c1457cc9145e13e936d90b3d9c7786b8b26cf4c7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{303, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2d051f91c5a9d440c5676985710483bc4f1a6c611b10c95a2ff0363d90c2a458, 256'h6ddf94e6fba5be586833d0c53cf216ad3948f37953c26c1cf4968e9a9e8243dc},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{306, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h530a0832b691da0b5619a0b11de6877f3c0971baaa68ed122758c29caaf46b72, 256'h6c89e44f5eb33060ea4b46318c39138eaedec72de42ba576579a6a4690e339f3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{309, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5924873209593135a4c3da7bb381227f8a4b6aa9f34fe5bb7f8fbc131a039ffe, 256'h1f1bb11b441c8feaa40f44213d9a405ed792d59fb49d5bcdd9a4285ae5693022},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{313, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h07dc2478d43c1232a4595608c64426c35510051a631ae6a5a6eb1161e57e42e1, 256'h4a59ea0fdb72d12165cea3bf1ca86ba97517bd188db3dbd21a5a157850021984},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{318, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2557d64a7aee2e0931c012e4fea1cd3a2c334edae68cdeb7158caf21b68e5a24, 256'h7f06cdbb6a90023a973882ed97b080fe6b05af3ec93db6f1a4399a69edf7670d},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{323, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5d5b38bd37ad498b2227a633268a8cca879a5c7c94a4e416bd0a614d09e606d2, 256'h12b8d664ea9991062ecbb834e58400e25c46007af84f6007d7f1685443269afe},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{324, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0c1cd9fe4034f086a2b52d65b9d3834d72aebe7f33dfe8f976da82648177d8e3, 256'h13105782e3d0cfe85c2778dec1a848b27ac0ae071aa6da341a9553a946b41e59},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{326, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h00a134b5c6ccbcefd4c882b945baeb4933444172795fa6796aae149067547098, 256'h566e46105d24d890151e3eea3ebf88f5b92b3f5ec93a217765a6dcbd94f2c55b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{327, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2e4721363ad3992c139e5a1c26395d2c2d777824aa24fde075e0d7381171309d, 256'h740f7c494418e1300dd4512f782a58800bff6a7abdfdd20fbbd4f05515ca1a4f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{328, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6852e9d3cd9fe373c2d504877967d365ab1456707b6817a042864694e1960ccf, 256'h064b27ea142b30887b84c86adccb2fa39a6911ad21fc7e819f593be52bc4f3bd},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{329, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h188a8c5648dc79eace158cf886c62b5468f05fd95f03a7635c5b4c31f09af4c5, 256'h36361a0b571a00c6cd5e686ccbfcfa703c4f97e48938346d0c103fdc76dc5867},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{331, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h07244865b72ff37e62e3146f0dc14682badd7197799135f0b00ade7671742bfe, 256'h0d80c2238edb4e4a7a86a8c57ca9af1711f406f7f5da0299aa04e2932d960754},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{334, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0bf6c0188dc9571cd0e21eecac5fbb19d2434988e9cc10244593ef3a98099f69, 256'h4864a562661f9221ec88e3dd0bc2f6e27ac128c30cc1a80f79ec670a22b042ee},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{336, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1cf3517ba3bf2ab8b9ead4ebb6e866cb88a1deacb6a785d3b63b483ca02ac495, 256'h249a798b73606f55f5f1c70de67cb1a0cff95d7dc50b3a617df861bad3c6b1c9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{338, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5f9d7d7c870d085fc1d49fff69e4a275812800d2cf8973e7325866cb40fa2b6f, 256'h6d1f5491d9f717a597a15fd540406486d76a44697b3f0d9d6dcef6669f8a0a56},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{339, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0a7d5b1959f71df9f817146ee49bd5c89b431e7993e2fdecab6858957da685ae, 256'h0f8aad2d254690bdc13f34a4fec44a02fd745a422df05ccbb54635a8b86b9609},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{340, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h79e88bf576b74bc07ca142395fda28f03d3d5e640b0b4ff0752c6d94cd553408, 256'h32cea05bd2d706c8f6036a507e2ab7766004f0904e2e5c5862749c0073245d6a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{342, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2664f1ffa982fedbcc7cab1b8bc6e2cb420218d2a6077ad08e591ba9feab33bd, 256'h49f5c7cb515e83872a3d41b4cdb85f242ad9d61a5bfc01debfbb52c6c84ba728},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{343, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5827518344844fd6a7de73cbb0a6befdea7b13d2dee4475317f0f18ffc81524b, 256'h4f5ccb4e0b488b5a5d760aacddb2d791970fe43da61eb30e2e90208a817e46db},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{345, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h52c683144e44119ae2013749d4964ef67509278f6d38ba869adcfa69970e123d, 256'h3479910167408f45bda420a626ec9c4ec711c1274be092198b4187c018b562ca},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{346, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h07310f90a9eae149a08402f54194a0f7b4ac427bf8d9bd6c7681071dc47dc362, 256'h26a6d37ac46d61fd600c0bf1bff87689ed117dda6b0e59318ae010a197a26ca0, 136'h014551231950b75fc4402da1722fc9baeb, 8'h03},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=136b(17B), s=8b(1B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h44ad339afbc21e9abf7b602a5ca535ea378135b6d10d81310bdd8293d1df3252, 264'h00b63ff7d0774770f8fe1d1722fa83acd02f434e4fc110a0cc8f6dddd37d56c463, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3e9a7582886089c62fb840cf3b83061cd1cff3ae4341808bb5bdee6191174177},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1260c2122c9e244e1af5151bede0c3ae23b54d7c596881d3eebad21f37dd878c, 256'h5c9a0c1a9ade76737a8811bd6a7f9287c978ee396aa89c11e47229d2ccb552f0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h24238e70b431b1a64efdf9032669939d4b77f249503fc6905feb7540dea3e6d2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1877045be25d34a1d0600f9d5c00d0645a2a54379b6ceefad2e6bf5c2a3352ce, 264'h00821a532cc1751ee1d36d41c3d6ab4e9b143e44ec46d73478ea6a79a5c0e54159, 8'h01, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h455439fcc3d2deeceddeaece60e7bd17304f36ebb602adf5a22e0b8f1db46a50, 264'h00aec38fb2baf221e9a8d1887c7bf6222dd1834634e77263315af6d23609d04f77, 8'h01, 8'h02},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2e1f466b024c0c3ace2437de09127fed04b706f94b19a21bb1c2acf35cece718, 256'h0449ae3523d72534e964972cfd3b38af0bddd9619e5af223e4d1a40f34cf9f1d, 8'h01, 8'h03},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008e7abdbbd18de7452374c1879a1c3b01d13261e7d4571c3b47a1c76c55a23373, 256'h26ed897cd517a4f5349db809780f6d2f2b9f6299d8b5a89077f1119a718fd7b3, 8'h02, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h7b333d4340d3d718dd3e6aff7de7bbf8b72bfd616c8420056052842376b9af19, 256'h42117c5afeac755d6f376fc6329a7d76051b87123a4a5d0bc4a539380f03de7b, 8'h02, 8'h02},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d30ca4a0ddb6616c851d30ced682c40f83c62758a1f2759988d6763a88f1c0e5, 256'h03a80d5415650d41239784e8e2fb1235e9fe991d112ebb81186cbf0da2de3aff, 8'h02, 8'h03},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{358, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h48969b39991297b332a652d3ee6e01e909b39904e71fa2354a7830c7750baf24, 264'h00b4012d1b830d199ccb1fc972b32bfded55f09cd62d257e5e844e27e57a1594ec, 8'h02, 24'hed2979},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=24b(3B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h02ef4d6d6cfd5a94f1d7784226e3e2a6c0a436c55839619f38fb4472b5f9ee77, 256'h7eb4acd4eebda5cd72875ffd2a2f26229c2dc6b46500919a432c86739f3ae866, 16'h0101, 256'h3a74e9d3a74e9d3a74e9d3a74e9d3a749f8ab3732a0a89604a09bce5b2916da4},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=16b(2B), s=256b(32B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h464f4ff715729cae5072ca3bd801d3195b67aec65e9b01aad20a2943dcbcb584, 264'h00b1afd29d31a39a11d570aa1597439b3b2d1971bf2f1abf15432d0207b10d1d08, 56'h2d9b4d347952cc, 256'h0343aefc2f25d98b882e86eb9e30d55a6eb508b516510b34024ae4b6362330b3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=56b(7B), s=256b(32B)
  '{361, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h157f8fddf373eb5f49cfcf10d8b853cf91cbcd7d665c3522ba7dd738ddb79a4c, 264'h00deadf1a5c448ea3c9f4191a8999abfcc757ac6d64567ef072c47fec613443b8f, 104'h1033e67e37b32b445580bf4efc, 256'h6f906f906f906f906f906f906f906f8fe1cab5eefdb214061dce3b22789f1d6f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=104b(13B), s=256b(32B)
  '{362, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0934a537466c07430e2c48feb990bb19fb78cecc9cee424ea4d130291aa237f0, 264'h00d4f92d23b462804b5b68c52558c01c9996dbf727fccabbeedb9621a400535afa, 16'h0101, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=16b(2B), s=256b(32B)
  '{363, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d6ef20be66c893f741a9bf90d9b74675d1c2a31296397acb3ef174fd0b300c65, 256'h4a0c95478ca00399162d7f0f2dc89efdc2b28a30fbabe285857295a4b0c4e265, 104'h062522bbd3ecbe7c39e93e7c26, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=104b(13B), s=256b(32B)
  '{365, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6e28303305d642ccb923b722ea86b2a0bc8e3735ecb26e849b19c9f76b2fdbb8, 256'h186e80d64d8cab164f5238f5318461bf89d4d96ee6544c816c7566947774e0f6, 72'h009c44febf31c3594d, 72'h00839ed28247c2b06b},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=72b(9B), s=72b(9B)
  '{366, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h375bda93f6af92fb5f8f4b1b5f0534e3bafab34cb7ad9fb9d0b722e4a5c302a9, 264'h00a00b9f387a5a396097aa2162fc5bbcf4a5263372f681c94da51e9799120990fd, 104'h09df8b682430beef6f5fd7c7cf, 104'h0fd0a62e13778f4222a0d61c8a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=104b(13B), s=104b(13B)
  '{367, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d75b68216babe03ae257e94b4e3bf1c52f44e3df266d1524ff8c5ea69da73197, 264'h00da4bff9ed1c53f44917a67d7b978598e89df359e3d5913eaea24f3ae259abc44, 136'h008a598e563a89f526c32ebec8de26367a, 136'h0084f633e2042630e99dd0f1e16f7a04bf},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=136b(17B), s=136b(17B)
  '{368, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h78bcda140aed23d430cb23c3dc0d01f423db134ee94a3a8cb483f2deac2ac653, 256'h118114f6f33045d4e9ed9107085007bfbddf8f58fe7a1a2445d66a990045476e, 168'h00aa6eeb5823f7fa31b466bb473797f0d0314c0bdf, 168'h00e2977c479e6d25703cebbc6bd561938cc9d1bfb9},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=168b(21B), s=168b(21B)
  '{369, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00bb79f61857f743bfa1b6e7111ce4094377256969e4e15159123d9548acc3be6c, 256'h1f9d9f8860dcffd3eb36dd6c31ff2e7226c2009c4c94d8d7d2b5686bf7abd677, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h01},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{370, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00bb79f61857f743bfa1b6e7111ce4094377256969e4e15159123d9548acc3be6c, 256'h1f9d9f8860dcffd3eb36dd6c31ff2e7226c2009c4c94d8d7d2b5686bf7abd677, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h00},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=8b(1B)
  '{371, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0093591827d9e6713b4e9faea62c72b28dfefa68e0c05160b5d6aae88fd2e36c36, 256'h073f5545ad5af410af26afff68654cf72d45e493489311203247347a890f4518, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h419d981c515af8cc82545aac0c85e9e308fbb2eab6acd7ed497e0b4145a18fd9},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{372, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h31ed3081aefe001eb6402069ee2ccc1862937b85995144dba9503943587bf0da, 264'h00da01b8cc4df34f5ab3b1a359615208946e5ee35f98ee775b8ccecd86ccc1650f, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h1b21717ad71d23bbac60a9ad0baf75b063c9fdf52a00ebf99d022172910993c9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{373, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h7dff66fa98509ff3e2e51045f4390523dccda43a3bc2885e58c248090990eea8, 256'h54c76c2b9adeb6bb571823e07fd7c65c8639cf9d905260064c8e7675ce6d98b4, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h2f588f66018f3dd14db3e28e77996487e32486b521ed8e5a20f06591951777e9},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{374, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4280509aab64edfc0b4a2967e4cbce849cb544e4a77313c8e6ece579fbd7420a, 256'h2e89fe5cc1927d554e6a3bb14033ea7c922cd75cba2c7415fdab52f20b1860f1, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h091a08870ff4daf9123b30c20e8c4fc8505758dcf4074fcaff2170c9bfcf74f4},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{375, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4f8df145194e3c4fc3eea26d43ce75b402d6b17472ddcbb254b8a79b0bf3d9cb, 256'h2aa20d82844cb266344e71ca78f2ad27a75a09e5bc0fa57e4efd9d465a0888db, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h7c370dc0ce8c59a8b273cba44a7c1191fc3186dc03cab96b0567312df0d0b250},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{376, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h009598a57dd67ec3e16b587a338aa3a10a3a3913b41a3af32e3ed3ff01358c6b14, 256'h122819edf8074bbc521f7d4cdce82fef7a516706affba1d93d9dea9ccae1a207, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h70b59a7d1ee77a2f9e0491c2a7cfcd0ed04df4a35192f6132dcc668c79a6160e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{377, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h009171fec3ca20806bc084f12f0760911b60990bd80e5b2a71ca03a048b20f837e, 256'h634fd17863761b2958d2be4e149f8d3d7abbdc18be03f451ab6c17fa0a1f8330, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h2736d76e412246e097148e2bf62915614eb7c428913a58eb5e9cd4674a9423de},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{378, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h777c8930b6e1d271100fe68ce93f163fa37612c5fff67f4a62fc3bafaf3d17a9, 264'h00ed73d86f60a51b5ed91353a3b054edc0aa92c9ebcbd0b75d188fdc882791d68d, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h4a1e12831fbe93627b02d6e7f24bccdd6ef4b2d0f46739eaf3b1eaf0ca117770},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{379, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00eabc248f626e0a63e1eb81c43d461a39a1dba881eb6ee2152b07c32d71bcf470, 256'h0603caa8b9d33db13af44c6efbec8a198ed6124ac9eb17eaafd2824a545ec000, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h06c778d4dfff7dee06ed88bc4e0ed34fc553aad67caf796f2a1c6487c1b2e877},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{380, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h009f7a13ada158a55f9ddf1a45f044f073d9b80030efdcfc9f9f58418fbceaf001, 264'h00f8ada0175090f80d47227d6713b6740f9a0091d88a837d0a1cd77b58a8f28d73, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h4de459ef9159afa057feb3ec40fef01c45b809f4ab296ea48c206d4249a2b451},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{381, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h11c4f3e461cd019b5c06ea0cea4c4090c3cc3e3c5d9f3c6d65b436826da9b4db, 264'h00bbeb7a77e4cbfda207097c43423705f72c80476da3dac40a483b0ab0f2ead1cb, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h745d294978007302033502e1acc48b63ae6500be43adbea1b258d6b423dbb416},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{382, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00e2e18682d53123aa01a6c5d00b0c623d671b462ea80bddd65227fd5105988aa4, 256'h161907b3fd25044a949ea41c8e2ea8459dc6f1654856b8b61b31543bb1b45bdb, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h7b2a785e3896f59b2d69da57648e80ad3c133a750a2847fd2098ccd902042b6c},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{383, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0090f8d4ca73de08a6564aaf005247b6f0ffe978504dce52605f46b7c3e56197da, 264'h00fadbe528eb70d9ee7ea0e70702db54f721514c7b8604ac2cb214f1decb7e383d, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h71ae94a72ca896875e7aa4a4c3d29afdb4b35b6996273e63c47ac519256c5eb1},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{384, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00824c195c73cffdf038d101bce1687b5c3b6146f395c885976f7753b2376b948e, 256'h3cdefa6fc347d13e4dcbc63a0b03a165180cd2be1431a0cf74ce1ea25082d2bc, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h0fa527fa7343c0bc9ec35a6278bfbff4d83301b154fc4bd14aee7eb93445b5f9},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{385, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2788a52f078eb3f202c4fa73e0d3386faf3df6be856003636f599922d4f5268f, 256'h30b4f207c919bbdf5e67a8be4265a8174754b3aba8f16e575b77ff4d5a7eb64f, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h6539c0adadd0525ff42622164ce9314348bd0863b4c80e936b23ca0414264671},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{386, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d533b789a4af890fa7a82a1fae58c404f9a62a50b49adafab349c513b4150874, 256'h01b4171b803e76b34a9861e10f7bc289a066fd01bd29f84c987a10a5fb18c2d4, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{387, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3a3150798c8af69d1e6e981f3a45402ba1d732f4be8330c5164f49e10ec555b4, 256'h221bd842bc5e4d97eff37165f60e3998a424d72a450cf95ea477c78287d0343a, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{388, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3b37df5fb347c69a0f17d85c0c7ca83736883a825e13143d0fcfc8101e851e80, 256'h0de3c090b6ca21ba543517330c04b12f948c6badf14a63abffdf4ef8c7537026, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a1},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{389, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00feb5163b0ece30ff3e03c7d55c4380fa2fa81ee2c0354942ff6f08c99d0cd82c, 264'h00e87de05ee1bda089d3e4e248fa0f721102acfffdf50e654be281433999df897e, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h44a5ad0bd0636d9e12bc9e0a6bdd5e1bba77f523842193b3b82e448e05d5f11e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{390, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h238ced001cf22b8853e02edc89cbeca5050ba7e042a7a77f9382cd4149228976, 256'h40683d3094643840f295890aa4c18aa39b41d77dd0fb3bb2700e4f9ec284ffc2, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h44a5ad0bd0636d9e12bc9e0a6bdd5e1bba77f523842193b3b82e448e05d5f11e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{391, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00961cf64817c06c0e51b3c2736c922fde18bd8c4906fcd7f5ef66c4678508f35e, 264'h00d2c5d18168cfbe70f2f123bd7419232bb92dd69113e2941061889481c5a027bf, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{392, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h13681eae168cd4ea7cf2e2a45d052742d10a9f64e796867dbdcb829fe0b10288, 256'h16528760d177376c09df79de39557c329cc1753517acffe8fa2ec298026b8384, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{393, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5aa7abfdb6b4086d543325e5d79c6e95ce42f866d2bb84909633a04bb1aa31c2, 264'h0091c80088794905e1da33336d874e2f91ccf45cc59185bede5dd6f3f7acaae18b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h16e1e459457679df5b9434ae23f474b3e8d2a70bd6b5dbe692ba16da01f1fb0a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{394, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 248'h277791b305a45b2b39590b2f05d3392a6c8182cef4eb540120e0f5c206c3e4, 256'h64108233fb0b8c3ac892d79ef8e0fbf92ed133addb4554270132584dc52eef41, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h1c940f313f92647be257eccd7ed08b0baef3f0478f25871b53635302c5f6314a},  // lens: hash=256b(32B), x=248b(31B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{395, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6efa092b68de9460f0bcc919005a5f6e80e19de98968be3cd2c770a9949bfb1a, 264'h00c75e6e5087d6550d5f9beb1e79e5029307bc255235e2d5dc99241ac3ab886c49, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h15d94a85077b493f91cb7101ec63e1b01be58b594e855f45050a8c14062d689b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{396, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h72d4a19c4f9d2cf5848ea40445b70d4696b5f02d632c0c654cc7d7eeb0c6d058, 264'h00e8c4cd9943e459174c7ac01fa742198e47e6c19a6bdb0c4f6c237831c1b3f942, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5b1d27a7694c146244a5ad0bd0636d9d9ef3b9fb58385418d9c982105077d1b7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{397, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2a8ea2f50dcced0c217575bdfa7cd47d1c6f100041ec0e35512794c1be7e7402, 256'h58f8c17122ed303fda7143eb58bede70295b653266013b0b0ebd3f053137f6ec, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2d85896b3eb9dbb5a52f42f9c9261ed3fc46644ec65f06ade3fd78f257e43432},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{398, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0088de689ce9af1e94be6a2089c8a8b1253ffdbb6c8e9c86249ba220001a4ad3b8, 256'h0c4998e54842f413b9edb1825acbb6335e81e4d184b2b01c8bebdc85d1f28946, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5b0b12d67d73b76b4a5e85f3924c3da7f88cc89d8cbe0d5bc7faf1e4afc86864},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{399, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00fea2d31f70f90d5fb3e00e186ac42ab3c1615cee714e0b4e1131b3d4d8225bf7, 264'h00b037a18df2ac15343f30f74067ddf29e817d5f77f8dce05714da59c094f0cda9, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h694c146244a5ad0bd0636d9e12bc9e09e60e68b90d0b5e6c5dddd0cb694d8799},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{400, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h7258911e3d423349166479dbe0b8341af7fbd03d0a7e10edccb36b6ceea5a3db, 256'h17ac2b8992791128fa3b96dc2fbd4ca3bfa782ef2832fc6656943db18e7346b0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3d7f487c07bfc5f30846938a3dcef696444707cf9677254a92b06c63ab867d22},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{401, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4f28461dea64474d6bb34d1499c97d37b9e95633df1ceeeaacd45016c98b3914, 264'h00c8818810b8cc06ddb40e8a1261c528faa589455d5a6df93b77bc5e0e493c7470, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6c7648fc0fbf8a06adb8b839f97b4ff7a800f11b1e37c593b261394599792ba4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{402, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h74f2a814fb5d8eca91a69b5e60712732b3937de32829be974ed7b68c5c2f5d66, 264'h00eff0f07c56f987a657f42196205f588c0f1d96fd8a63a5f238b48f478788fe3b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h641c9c5d790dc09cdd3dfabb62cdf453e69747a7e3d7aa1a714189ef53171a99},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{403, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h195b51a7cc4a21b8274a70a90de779814c3c8ca358328208c09a29f336b82d6a, 264'h00b2416b7c92fffdc29c3b1282dd2a77a4d04df7f7452047393d849989c5cee9ad, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h29798c5c45bdf58b4a7b2fdc2c46ab4af1218c7eeb9f0f27a88f1267674de3b0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{404, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h622fc74732034bec2ddf3bc16d34b3d1f7a327dd2a8c19bab4bb4fe3a24b58aa, 256'h736b2f2fae76f4dfaecc9096333b01328d51eb3fda9c9227e90d0b449983c4f0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h0b70f22ca2bb3cefadca1a5711fa3a59f4695385eb5aedf3495d0b6d00f8fd85},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{405, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1f7f85caf2d7550e7af9b65023ebb4dce3450311692309db269969b834b611c7, 256'h0827f45b78020ecbbaf484fdd5bfaae6870f1184c21581baf6ef82bd7b530f93, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h16e1e459457679df5b9434ae23f474b3e8d2a70bd6b5dbe692ba16da01f1fb0a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{406, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h49c197dc80ad1da47a4342b93893e8e1fb0bb94fc33a83e783c00b24c781377a, 264'h00efc20da92bac762951f72474becc734d4cc22ba81b895e282fdac4df7af0f37d, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2252d685e831b6cf095e4f0535eeaf0ddd3bfa91c210c9d9dc17224702eaf88f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{407, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d8cb68517b616a56400aa3868635e54b6f699598a2f6167757654980baf6acbe, 256'h7ec8cf449c849aa03461a30efada41453c57c6e6fbc93bbc6fa49ada6dc0555c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h75135abd7c425b60371a477f09ce0f274f64a8c6b061a07b5d63e93c65046c53},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{408, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h030713fb63f2aa6fe2cadf1b20efc259c77445dafa87dac398b84065ca347df3, 264'h00b227818de1a39b589cb071d83e5317cccdc2338e51e312fe31d8dc34a4801750, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa3e3a49a23a6d8abe95461f8445676b17},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{409, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00babb3677b0955802d8e929a41355640eaf1ea1353f8a771331c4946e3480afa7, 256'h252f196c87ed3d2a59d3b1b559137fed0013fecefc19fb5a92682b9bca51b950, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3e888377ac6c71ac9dec3fdb9b56c9feaf0cfaca9f827fc5eb65fc3eac811210},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{410, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1aab2018793471111a8a0e9b143fde02fc95920796d3a63de329b424396fba60, 264'h00bbe4130705174792441b318d3aa31dfe8577821e9b446ec573d272e036c4ebe9, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h30bbb794db588363b40679f6c182a50d3ce9679acdd3ffbe36d7813dacbdc818},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{411, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008cb0b909499c83ea806cd885b1dd467a0119f06a88a0276eb0cfda274535a8ff, 256'h47b5428833bc3f2c8bf9d9041158cf33718a69961cd01729bc0011d1e586ab75, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2c37fd995622c4fb7fffffffffffffffc7cee745110cb45ab558ed7c90c15a2f},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{412, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008f03cf1a42272bb1532723093f72e6feeac85e1700e9fbe9a6a2dd642d74bf5d, 256'h3b89a7189dad8cf75fc22f6f158aa27f9c2ca00daca785be3358f2bda3862ca0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h7fd995622c4fb7ffffffffffffffffff5d883ffab5b32652ccdcaa290fccb97d},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{413, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h44de3b9c7a57a8c9e820952753421e7d987bb3d79f71f013805c897e018f8ace, 264'h00a2460758c8f98d3fdce121a943659e372c326fff2e5fc2ae7fa3f79daae13c12, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 248'h4cd53ba7608fffffffffffffffffffff9e5cf143e2539626190a3ab09cce47},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=248b(31B)
  '{414, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6fb8b2b48e33031268ad6a517484dc8839ea90f6669ea0c7ac3233e2ac31394a, 256'h0ac8bbe7f73c2ff4df9978727ac1dfc2fd58647d20f31f99105316b64671f204, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5622c4fb7fffffffffffffffffffffff928a8f1c7ac7bec1808b9f61c01ec327},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{415, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00bea71122a048693e905ff602b3cf9dd18af69b9fc9d8431d2b1dd26b942c95e6, 264'h00f43c7b8b95eb62082c12db9dbda7fe38e45cbe4a4886907fb81bdb0c5ea9246c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h44104104104104104104104104104103b87853fd3b7d3f8e175125b4382f25ed},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{416, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00da918c731ba06a20cb94ef33b778e981a404a305f1941fe33666b45b03353156, 264'h00e2bb2694f575b45183be78e5c9b5210bf3bf488fd4c8294516d89572ca4f5391, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2739ce739ce739ce739ce739ce739ce705560298d1f2f08dc419ac273a5b54d9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{417, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3007e92c3937dade7964dfa35b0eff031f7eb02aed0a0314411106cdeb70fe3d, 256'h5a7546fc0552997b20e3d6f413e75e2cb66e116322697114b79bac734bfc4dc5, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h4888888888888888888888888888888831c83ae82ebe0898776b4c69d11f88de},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{418, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h60e734ef5624d3cbf0ddd375011bd663d6d6aebc644eb599fdf98dbdcd18ce9b, 264'h00d2d90b3ac31f139af832cccf6ccbbb2c6ea11fa97370dc9906da474d7d8a7567, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6492492492492492492492492492492406dd3a19b8d5fb875235963c593bd2d3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{419, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0085a900e97858f693c0b7dfa261e380dad6ea046d1f65ddeeedd5f7d8af0ba337, 256'h69744d15add4f6c0bc3b0da2aec93b34cb8c65f9340ddf74e7b0009eeeccce3c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa3e3a49a23a6d8abe95461f8445676b15},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{420, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h38066f75d88efc4c93de36f49e037b234cc18b1de5608750a62cab0345401046, 264'h00a3e84bed8cfcb819ef4d550444f2ce4b651766b69e2e2901f88836ff90034fed, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa3e3a49a23a6d8abe95461f8445676b17},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{421, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0098f68177dc95c1b4cbfa5245488ca523a7d5629470d035d621a443c72f39aabf, 264'h00a33d29546fa1c648f2c7d5ccf70cf1ce4ab79b5db1ac059dbecd068dbdff1b89, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffe},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{422, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5c2bbfa23c9b9ad07f038aa89b4930bf267d9401e4255de9e8da0a5078ec8277, 264'h00e3e882a31d5e6a379e0793983ccded39b95c4353ab2ff01ea5369ba47b0c3191, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h185ddbca6dac41b1da033cfb60c152869e74b3cd66e9ffdf1b6bc09ed65ee40c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{423, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2ea7133432339c69d27f9b267281bd2ddd5f19d6338d400a05cd3647b157a385, 256'h3547808298448edb5e701ade84cd5fb1ac9567ba5e8fb68a6b933ec4b5cc84cc, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 256'h29ed3d67b3d505be95580d77d5b792b436881179b2b6b2e04c5fe592d38d82d9},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{424, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2ea7133432339c69d27f9b267281bd2ddd5f19d6338d400a05cd3647b157a385, 264'h00cab87f7d67bb7124a18fe5217b32a04e536a9845a1704975946cc13a4a337763, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 256'h29ed3d67b3d505be95580d77d5b792b436881179b2b6b2e04c5fe592d38d82d9},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{425, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008aa2c64fa9c6437563abfbcbd00b2048d48c18c152a2a6f49036de7647ebe82e, 256'h1ce64387995c68a060fa3bc0399b05cc06eec7d598f75041a4917e692b7f51ff, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0, 256'h33333333333333333333333333333332f222f8faefdb533f265d461c29a47373},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{432, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3f3952199774c7cf39b38b66cb1042a6260d8680803845e4d433adba3bb24818, 256'h5ea495b68cbc7ed4173ee63c9042dc502625c7eb7e21fb02ca9a9114e0a3a18d, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{433, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00cdfb8c0f422e144e137c2412c86c171f5fe3fa3f5bbb544e9076288f3ced786e, 256'h054fd0721b77c11c79beacb3c94211b0a19bda08652efeaf92513a3b0a163698, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{434, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h73598a6a1c68278fa6bfd0ce4064e68235bc1c0f6b20a928108be336730f87e3, 264'h00cbae612519b5032ecc85aed811271a95fe7939d5d3460140ba318f4d14aba31d, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{435, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h58debd9a7ee2c9d59132478a5440ae4d5d7ed437308369f92ea86c82183f10a1, 256'h6773e76f5edbf4da0e4f1bdffac0f57257e1dfa465842931309a24245fda6a5d, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{436, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008b904de47967340c5f8c3572a720924ef7578637feab1949acb241a5a6ac3f5b, 264'h00950904496f9824b1d63f3313bae21b89fae89afdfc811b5ece03fd5aa301864f, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{437, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f4892b6d525c771e035f2a252708f3784e48238604b4f94dc56eaa1e546d941a, 256'h346b1aa0bce68b1c50e5b52f509fb5522e5c25e028bc8f863402edb7bcad8b1b, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{439, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 256'h44a5ad0bd0636d9e12bc9e0a6bdd5e1bba77f523842193b3b82e448e05d5f11e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{441, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 256'h44a5ad0bd0636d9e12bc9e0a6bdd5e1bba77f523842193b3b82e448e05d5f11e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{443, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h109cd8ae0374358984a8249c0a843628f2835ffad1df1a9a69aa2fe72355545c, 256'h5390ff250ac4274e1cb25cd6ca6491f6b91281e32f5b264d87977aed4a94e77b},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{445, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h4f053f563ad34b74fd8c9934ce59e79c2eb8e6eca0fef5b323ca67d5ac7ed238, 256'h4d4b05daa0719e773d8617dce5631c5fd6f59c9bdc748e4b55c970040af01be5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{446, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h6d6a4f556ccce154e7fb9f19e76c3deca13d59cc2aeb4ecad968aab2ded45965, 256'h53b9fa74803ede0fc4441bf683d56c564d3e274e09ccf47390badd1471c05fb7},  // lens: hash=256b(32B), x=256b(32B), y=232b(29B), r=256b(32B), s=256b(32B)
  '{449, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h3854a3998aebdf2dbc28adac4181462ccac7873907ab7f212c42db0e69b56ed8, 256'h3ed3f6b8a388d02f3e4df9f2ae9c1bd2c3916a686460dffcd42909cd7f82058e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{451, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h49fc102a08ca47b60e0858cd0284d22cddd7233f94aaffbb2db1dd2cf08425e1, 256'h5b16fca5a12cdb39701697ad8e39ffd6bdec0024298afaa2326aea09200b14d6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{452, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h41efa7d3f05a0010675fcb918a45c693da4b348df21a59d6f9cd73e0d831d67a, 256'h4454ada693e5e26b7bd693236d340f80545c834577b6f73d378c7bcc534244da},  // lens: hash=256b(32B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{455, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'h62f48ef71ace27bf5a01834de1f7e3f948b9dce1ca1e911d5e13d3b104471d82, 256'h5ea8f33f0c778972c4582080deda9b341857dd64514f0849a05f6964c2e34022},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{458, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'h592c41e16517f12fcabd98267674f974b588e9f35d35406c1a7bb2ed1d19b7b8, 256'h3e65a06bd9f83caaeb7b00f2368d7e0dece6b12221269a9b5b765198f840a3a1},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{461, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h176a2557566ffa518b11226694eb9802ed2098bfe278e5570fe1d5d7af18a943, 256'h1291df6a0ed5fc0d15098e70bcf13a009284dfd0689d3bb4be6ceeb9be1487c4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{462, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h60be20c3dbc162dd34d26780621c104bbe5dace630171b2daef0d826409ee5c2, 256'h427f7e4d889d549170bda6a9409fb1cb8b0e763d13eea7bd97f64cf41dc6e497}  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
};
`endif // WYCHERPROOF_SECP256K1_SHA256_V1_SV
