`ifndef WYCHERPROOF_SECP224R1_SHA3512_SV
`define WYCHERPROOF_SECP224R1_SHA3512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224r1_sha3512;

localparam int TEST_VECTORS_SECP224R1_SHA3512_NUM = 79;

ecdsa_vector_secp224r1_sha3512 test_vectors_secp224r1_sha3512 [] = '{
  '{144, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{232, 1'b1, 512'h4a00000000d34b9c928306129f1a8059b199049f30ffd4d5b9747c848b197497634fb5190298af2f6a90d273164d68431c984e0fcd3a810ccd7b95b5e0dcd21f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1bb6ce51b7e504ccd69a910a11a9c29ba77100d5bccb179de19a93dd, 224'h770a160b2635bb293c73a07fb1fd5e0314b50127ab3e70d1ab974de6},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{240, 1'b1, 512'hb1fe8fe86f9994808c00000000f313a999ae7b5281bcacf933f05e4c8d526e761afa3141e9efefe959438620220c28bbad7047a6c1a98f95520baeb1d7af6278, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h398b59d0b6a7171d3518d1d3ef6796f10a14251aca5630fa32655741, 224'h4259d0edc9c2aabc09c37a69444df24a5191e21d387b98b080745279},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{242, 1'b1, 512'hed19e69c6f4de76b35ce6c00000000ad94175b8ad5f1fb69995d7d87abd893772b81ff83fd6caa25d1fe69b0317ec4068cdddac49512e6bf12d9cd8ce9a951c7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7f5127a83c76554fe4fcc00ea6e62b14c8a675168e60ea9d6b1f034d, 224'h7ab4aca6a9315c795936fb41bcf46a4840a1e41a874ddb1ad5b550a7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{249, 1'b1, 512'hd912418a7d72e83ab66eed185bd627c70b00000000a88db442365b3ec21269abd09b4b2e040304518850835236add11fecca5a2c529f8bc4c06174a03b997830, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b00ebcedc8c30521024d15dfa14304f8c594ab8a17eb3df68393b2e, 224'h3a53183103dd1b1ef8631e7cafe510eac9ab4c10164df208c598e20f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{251, 1'b1, 512'h91f07f1a3d4b600628f1754ae5ec28d43554a40000000051e8c4594c5a2e68bf2f497bfbc7e703e1b18398a0b5515a38d60284b1a2dfad8c9132a7b9a98db6eb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h504f2f50ca931e2a4f8cda0f08c2b79ef051677d76a08f1806c53af5, 224'h736248501f062b14bd3fee6528700d1a64a8ae30d7c76e1a92b66bad},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{253, 1'b1, 512'h7da7793b2bed3ce23ef7f1c04376791fa03f741f650000000008744fe10ac37fab4edf76492a339fe79e56ef75aee6c3169a0a61e3cb27e74666a4fe4184526c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h32377296ba47114b5f3dcff841416bca3e5e98d64dd987badc457655, 224'h29a37a143b47b029e256c7506a679ee8f1962ccbbb1c83f4088501b2},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{254, 1'b1, 512'h48cd33f55583315ab2131d5db1f9cfcb0590b13a266700000000c9bd5d6fbcdf457e3bffd7b4875145a47be68b99a201b93b8685e80d61ce692a913be1183569, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h75d62c172f26e6e6831c233b49895c1a87c1ee3ef57b711856199e46, 224'h27830a8d1fc44993990a9d1b2b147ff8792b0b0823bc30fb012ce9ee},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{257, 1'b1, 512'h90f9b7739bb1699b90bfdf7cef079649e3f08242a08d05026100000000d3a4568eccd5ef4d94de4885986b68670617f552b9cb2a6eed337392b49ad4d04a9dad, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1a71aa363800731f4c5a9f0a4235198a7658f1b425972ecac9a2a340, 224'h21b61939e575b1a5ff487473ba3803683c8b20e89844a55785630f89},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{263, 1'b1, 512'hdfe80a6b887fa09cbdc8bb94300a4ad38f0380331a18c0a0b62708e590dd3800000000d364091041bb72f35391e792802f5c23fd676d0775e56ac2e41880d92d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0fc1582e0b3ebe74b1fa4425e321a5b2d16b1c3ab060e98cf530defa, 224'h115eae025fa3422621a49fd78486ca245894a2d83c644e31abe21b5b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{295, 1'b1, 512'h9481ffffffff6e35dfab283e61e8f9a49de1cda44cdf1e2680292ded627b16d9b566ac057cef4c3380ee126c020a6ae86ded132faef613440c54185ed5986dcd, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h565c6827c8f18daa21a6b1edb8af81193e8e391f3e8360b346c7b98a, 224'h468b8b2e16c51e41e26651493e02f0db3af5c9981edfff2991d10599},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{296, 1'b1, 512'h2d8fbaffffffffb42e8498ddf2697ff4a2223fac0c486f05f57374d84dab9e8d13f52f6c898c8a7a74f2d48bee3cc16265e12a6dca3bee77c0ff0ee5e9af7e49, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6030ec07ae1cd991dfbc6b48da43c6240b5bb8f7fe19832df596754d, 224'h54b93d4ae52e4cb7eb969a1eb62f0be395d30a43e7d5736df6b508fc},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{301, 1'b1, 512'hc17991fc38743c0bffffffff12be8c0818873e8d65ea350547aa4cdc067cd0a4c21e1d9387ca3c60306f95160cc1f85a08ebdd4f3107b359483b719f5b9a18ab, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5dd7d39e95169cefd77a5a5dfd435e2a879576faf3a845d266d402ca, 224'h63225084b9219b15884e0cd665aca92ef1f4b541987b98cbd03edbfb},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{303, 1'b1, 512'he4d30dcc9e0b433fac32ffffffff83bb0169390c4443bfa7b7bc8a7c4421fb94a64d266b35ee622ee92a194a9c369a1bdd0961e4047a4fc3ed632b51f01547c1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h16881c4ae60f32a6b81d445f7bb921ce4f4dcd349695efe0fc94d213, 224'h06066332f61edc98a88a21a42f26e912c99c5471093aca9b1c11d54e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{304, 1'b1, 512'h8f46b06e493783b6d3209bffffffff5f263101ceb63bd0313945c63e59a123011230ea2a874c147574859882f49e6fdc842cbd97843daff440629f6a58573ee8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3d0af397602fc0d18d8a733377cc3e596c143f75d6a9d2c62c99f327, 224'h30ad8bf0bef3b8a2bb4158db621de4570d75c5fec7bb8c3e78af8445},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{312, 1'b1, 512'hffde6b2d174d86702f3a46946c7167cabd18feffffffff2df58cb555aad0b0df043b0c01b91bf2ee4827aac1d987f3174e1fce7921c831a0b0aeab1ad1156fed, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h32c28f726d79d4610f6382c329a3a955059f5876ef343585098f40db, 224'h20d7df0ae11f3909ffdc54b12d05bd294505ab76058c79c61dfceedd},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 512'hc0635b12b9164d0a9480ba133839afb60f79f6e7fa22fffffffff18d9363b5c503a5ae2f4cea06d8c5333965149a2cd0ed0491d1f9c8cfbf12fce9914dc22f30, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h431e666843a0d5e131567ab13ec0accd1fef8d441e96c4b8834d4e40, 224'h0e7a8bb3cef5a676cf4148da42b61457cf9fd43c8a33241d4bb87181},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{321, 1'b1, 512'hef503ce85b5b48ef35abff5d47345a71aa715f5e8e1568c9721a78ffffffffffe6124c567f2fb5b5f476271da455e079b655dc8c9506b65d9e3c60892984e8ba, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h762764cf2163759dfcf7863b20849c6deb57808cb208479814a243f8, 224'h7b41a973df219ea717a653bdbe27669bba57fc7c7afc3afe9c87d62f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{323, 1'b1, 512'h9e670958749c5bbc0cacb1ee6c38e71eede821d75d84cc2fe1335af9f6ffffffff4e9613cec31f535c4c7bdab269d70a8d4b3bdffa3065d91435a4237cae96da, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h531c06348905bbf16d85b8eba22f5d5ca33e490107ea979f6f322a65, 224'h0109215bf6d2afbedf4efe481f704963355f09f59e1977be330972a7},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{325, 1'b1, 512'h59f9626626a34d5491d567d0315894fb702c1d7a2ec677a2b595a772b20d8effffffff20557e965f33f606242a59aea4cd565aecb931664e51fee93a92ccaab6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70ba414a666f89e84064b2f9b08d500c6bb12d0a5ef9b23f4fa46ccf, 224'h43d88b7e943fe8792ff62ed462ea308d28f7f03e4dc59d6214f30507},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{335, 1'b1, 512'h4e29d13bd24e9f13d5e31ac769469a23d44278a67b110f7bab6095667a3a5180bc8124849e31af47ffffffff94e438c9abcb1301833210026c068417d2da4b20, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6808f8c1cf3a051724d074ebdc85fcdc14987324605a81db7591baa6, 224'h026f5efef2c657bc048c88a165f885628efcad293d80a5cf72855491},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{337, 1'b1, 512'h7692bad59be557b4e1db6cf148e5f0ff3c273d29d9017b90c8c26236cf78465b335a40716400ae0aaa34ffffffffd68ebefa85c403e0a25dbfeda3354bcc2a84, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4cb87503bde0aca323f93b04e1735f84bc0e101ba8b71332fb40ce4c, 224'h0bbc59dac149a5644771119b00d1d72905e4b080f9aff5d6a42e1565},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{343, 1'b1, 512'h388b354799942c6595ba49bc6bf8e7ca5c06c6ae8015c0f58e69192d96cc60e30696c1284ba98c1b22c5c7f23bf8e0ffffffff15f579e355c7258262f0fdfdfb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h733752fa2b90121c01878170f2019d9c9a4b1c95e82acab18ae95d71, 224'h358eb5d69942b4b5d0d900bb843d79f90af54663b3a926fabd081d42},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{344, 1'b1, 512'hc6bf307fea8c2799ef482911ac86779072e5757f934a3671ad8c5a9e372bb2ec8d318ee3bd0cc4460f9050c937a3409cffffffff81c81c22e9468fd07ec09f55, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h72fa0cb38863c06e535402e010bac709ef4beb0b38118c7b13308e83, 224'h33eb21f6c081afa7db62c2f8cf78ed1982cb762a130509bdb53f1774},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{346, 1'b1, 512'hd88d68932ee321d611334d87de84ef4240025f9d0c8f11bd9aaea2e7729ad87ab0ee66d229b2eb78221050b375a54bd698a2ffffffff0967dbcb983a8f09417c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h37e05ebb376ede0d3fc7528f19dbe4a38e4f310295058e2173f88900, 224'h4f8d5ca627d43c54db6674e1462d12c42603cddc6f3067307ab04d4f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{348, 1'b1, 512'h4f34828f9520f17da9e588884a26df5ab85e8456184bb19001abc926a180c32a112ba4164e81d69b8fdaaf3c60619a7d1a5840b6ffffffff8748db5ab09c4a64, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h05ea0f04e9b4eb3b62fcf8f1f1d120e58a932ca9a04e8c64bbee537e, 224'h166633a3c8d2b5c6246da69e069f2f09a7912efc355c405302b2984b},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{351, 1'b1, 512'h0844602883dbcf60972c8b943b5ea020ccb0d19c82eb86cb18d4225a79f97279539214d6e3df6ba6af165c9cd95b8b67a36b39bbd101ffffffff5a9aa9794dd2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1bc64aaf83515275fd3187a18d3651c75ce85b53f5579ecf5f190334, 224'h2ed9fc723bd723cd4c8b62b7968e5f058d25aa6f6bb45e6b09337793},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{352, 1'b1, 512'h73672c1037e14e2ed10a0928e8938944667e83879d16f2688f2fe0087494b9f496471dd4e27f5cfddfc4b5efc4e7fcd511d2f67ea879f2ffffffffaebc4501e4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h240d8b05889274d716f57588536320775afed824d79f41f32c35e728, 224'h25031a073d638165f8c0b46a28e008f1de9fa0cf726d316269f669d6},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{362, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h448bad17b638f55372b256c6717ac0fe443c20af133348be8f728577, 224'h421c701ae6015da98a2ec4140122091588c013a74fd78b3814c981b2, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{364, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00fad98df6a5fbd9f3c023f2ab809c57c72de3396d1cae4bc35d78d8d1, 232'h00889e372a90189ece8fbc690fe3cdeeef38ab12ffda721f32f849ae50, 8'h03, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{365, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00d2eaeb6be6b5dced48d595b95f73b069f49a078572c74dbc557fa25a, 232'h00a6388c4362e6aa12ab9c1350cd6789d0955445d9198ecc3a4618da73, 8'h03, 8'h03},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{366, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h2df6ce6019d77e3c6e04908a3fde5b8833f9c493bf3cc6568e3d40cb, 224'h0ced2e9cad2ed363fd20aeb9983bcb22091fcb559c1f6fd538a0ae04, 8'h03, 8'h04},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{370, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h008f711e9fbea41bd25aadf584999926a29c2801e7dbb2eb1dbe0d1586, 232'h00841a143bdeeac9969be87f57b4d71a466b2b6aed24e854b07570e629, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=56b(7B), s=224b(28B)
  '{371, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00c288ddd81714a9e766b35a03c835fbe1a52c540b747b11ba3ebabdcc, 232'h00b26bd049bd3088b553162261eb93ab5a75d873bfca8122a229e2cfc7, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{375, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00c847d6757702db5d47caf6129e865aa22d6b55c545f70ce7e7ad0eca, 232'h00f69bf4c624111ef1ce92e9e10d126f0ceda9851dcc53993930324d3e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{376, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00c847d6757702db5d47caf6129e865aa22d6b55c545f70ce7e7ad0eca, 232'h00f69bf4c624111ef1ce92e9e10d126f0ceda9851dcc53993930324d3e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{377, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h61c0d09fc40dd59a7b5281af54fd4db8819997cf31212a4b35cf6078, 232'h00a55ef14cafacd57ca50195aa1962aa7d01f7595d76d342d83fed44ec, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{378, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h66539275c7d5ae5dad2507a7169c48a9cff067c4d6afeb22561239b6, 224'h12eec9a7e63d602cf87f3581bdeb19ce994c48b41079ef8186339dfd, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{379, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h43a45adf3cd2a866e01ec45269f604af026a4483973cc4356b473966, 224'h2a8403f5f14fcd737d2aedec136a534417e0d19e1b98d53944100d0f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{380, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h2e55f92435ee396708e4805e3a2c4c6152c69e1671e9d6387c56f58d, 224'h3b4a173ad9f475448586ae0f531ee07f15553eba9828b2bc8d72c5f1, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd543},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{382, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h144765b9d78724babc4358b229df98e9d64da22724381ebfe41d7e72, 232'h0086e958c2f6779b8ea76433cd4dce0ae4cd300875ac1c7ad218e57a55, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{385, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00d2612ed20fe786484b8955d658200776ec219426479c69194f8c1baf, 232'h00a3af3aa778c1751f4474cc0ff2db2a834c232ec49e9ce142a51170b7, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2d4465a55b282f252f2b47f9f7bfc0ba40ec4dca29f567940b2d90f4},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{386, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h4c70cd0aa06d9ee36a16202bcfc891ceb41a26e0bcdde9d93da8001a, 232'h00ab77b507c77931fc7ee290cda7b7af6ad90d0c97b836ae1b65b6eccb, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fe808b87e0e6e76364ce32fde12f692d69dd3b362ef4cf499e03418},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{388, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h79e577f8303d4ed74c3a19cabe3ec35bd39cb789bc7309335a5710e6, 224'h43cc437d5793931f92eea56039b22088165693a7d9ed0ffc6188aa24, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c957342d757ecbd2518ae59c5c2f4ebdd95caedf61c68b89387f3c9},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{390, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00ee2558b8b7642287cdeedc8bca740974264a667e5edefe79e7a03900, 224'h5cf362e47faca649cf9b8f6c9214539ef2eee6b86935185c1fdb3492, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h342d757ecbd2518ae59c5c357e76013b79f087e62e58923f7ea5c045},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{391, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00f8b4c378bd5f417b562ae127f39825a2b05770089b7caf9324d7ce1a, 224'h50708175ba245e9c152bff3ca95743e261b6f579328f30680fb6a2a0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h21f862ec7b9a0f5e3fbe5d774e20a59eb3c341b9e1ff215b446f637f},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{392, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h5eb63f0f7b7ec667588670022e2f0b1124b132ebe16c143d6ed24602, 232'h00af2b27b92a449a4edc20267d25d0a238b43aa7289348a1378db079de, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h43f0c5d8f7341ebc7f7cbaee9c414b3d67868373c3fe42b688dec6fe},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{393, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h280ac7f11afa66465c37eba820aa8f393d13c5634022333c7a2524bd, 224'h5c63b1e9ed18115b589b56270c5c3281fa97060f1d30aef465f445e2, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h65e928c572ce2e1abf3b1865ea61f0dc1b49c52da5fd6411cd4e2a7d},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{394, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00cdc63e73d8d6f4f8770a97d93bde4e1974a277adad53d500cb070907, 224'h533c09379488cb344ce01bb29a2f12d6e0b946a279c7f5d47831477c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3ff4045c3f07373b1b267197ef097b496b4ee9d9b177a67a4cf01a0c},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{395, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h5e963ce90708539b001d821b9884f46ee4ba452bfcd539741d8fe838, 224'h4c8dc874329bd0b78fe04e0291f13907ff5723e8d15146c5469d7d9b, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{397, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b97529fb4a1e02b5e81d77b0e7909a2fde857a1edc9fa660d600c89a, 232'h00e5a8c9c55885cc20f54f5c8f423f785caf423d77ba0afc31fc16f131, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{399, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00d656048bfd65af83d6dc3f7cb7d240c9e0cdee6e946b15abb13f4b33, 232'h00d61580a159caf9fd87194b7c9d78753e0e00560a208d34c7dd4c6a63, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{401, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00912cff3ab4338f1f09b71f909dd68186cfabeb746beae33700dd923f, 232'h00f832461ccff9b83c25754bc1def8f10c5ffbdca0127914cf24184823, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{403, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h0086ec9d3ba7c6d9498069a07761a9d85e04fa21fd599c6a2664e86254, 232'h00c5900aa4b9882b32983c5e029fe6a5578ac818e79acb20beef73e8ee, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{404, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b08c34e9416743b6a3f52c42041a5fc3011f64dffb54875bc690393e, 224'h6a7c67833682e81719f928df55faac24f488028515b26e03c1c9a02c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{408, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b08c10bbd277ee6ab501aa71141733cb196b74de463ead5ea224022c, 224'h7f68bcdeead7d74cb6186e32219846424a926dec60b2a227411ae805, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{409, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b1babefd03f6f738fc86d32ca245f5db21f67e7bd919079bd735f35b, 232'h00d9ad5e6886dcfc7f2272b98c48a7c43f1c57a024f2f054fc59bb4354, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{411, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00f9973f688705dc1025beb72663df6f84bda4a14a79e5953d699269ba, 232'h00886f01e609345596494468378d758c618f49e216287d85554af8eb68, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{413, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h0ac469e816565a6a74bec821ca20b88a61018a0335199b5d7bd969e9, 224'h463355c73a2d9c51049f7a94509a9ac4ea0165763ba113a30db999e2, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=512b(64B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{414, 1'b1, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 224'h662eb328d24fb548f51792b5563ac3cb237f0a65199460eebfcaa5c3, 232'h00e758d13e7b419b417c8c97c4727c39fd373045e18792ad8076b072b4, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{421, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd543, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{423, 1'b0, 512'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd5435447f1c3a56f87db98089d208c89e902bb50ed289995ee7ccf6d6e6b1cec4aaf832d3734, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h342dae751a63a3ca8189cf342b3b34eaaa2565e2c7e26121c1bfd543, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{428, 1'b1, 512'h7d795fe6a97761d89b35f64e09555951f6ec2a669a9fa03481c100ae158f183e2171e142437d2c3a42352108a22a7e3d797beaf6c3075db419b6f4acca479c83, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h0316a2259370447c1b06f51f6189b033ead956c11ebbc3edbdc2b5e4, 224'h24bda2d065a0475c9fc5ee300f6c4c826b07a740d4990fcc146006aa},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{439, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h3fdb17cc44c9a0e995290a458c2f64b8565541cf56139575212ec168, 224'h5e51c778b560f3c61bc3bf0eb50ff8d34dcb5eb85cc25b4ae6a7443a},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{440, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h1d98253a63b83f0e042ed2c342fd4217c29f990fcd5b5cbb9e51721f, 224'h49fcf5e4d680cdd36405c514414cc47d9731a97c4edcbac7b7b27f89},  // lens: hash=512b(64B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{443, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h4d96e743ac0dbbf2413725a193c7e70947b59501601e337665023ee2, 224'h764ef71a184f0244c0e1de1b729b8421be53bd0ded2015dc3d1f1a13},  // lens: hash=512b(64B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{444, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h060ac961eff4e5053f7045b9ea1db338dd4b3a6cce331386d3988655, 224'h0cfc61a43a67d0660fc386efc1b603b28f651885bff519c632e11a8c},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{445, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h3415d0790d9b9ba8ffa82f447a4fed58cce3ebbaf43b68c162495c85, 224'h1e0e20ac93d19dbd9ddd632e5c0910560e941acf2ba5d7f3f2abe27f},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{446, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h2066593be10db4111e032cce79004a2e66aff1774d595ad4c37b61d6, 224'h2aaddfe2abcbb137ebf80d35c86c7f81fc760640eec39eb3abe9ee7d},  // lens: hash=512b(64B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{448, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h2d738785b04282261457a9b149a6c51c4c611f29e14113bbd2625981, 224'h6cacb7671751394b931ab86a09631ee26cd077c01af8c3491b535982},  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{449, 1'b1, 512'h740913294202f7597ef7c2ae48b64b02482e698abf5c4fbbc85c7c321e10bfb22050f90fba281c46f15a058697bb7e5112bdfcdbf656bc61bd7b3b2678b548a6, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h121f5992ff2892a8e0b36cf4f31331fddcb9b53d1aec2c7d9cd887cb, 224'h406a219f572c58baab779d8c386fe8e84857024a21c01f949505a668}  // lens: hash=512b(64B), x=200b(25B), y=232b(29B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224R1_SHA3512_SV
