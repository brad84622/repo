`ifndef WYCHERPROOF_SECP256K1_SHA512_SV
`define WYCHERPROOF_SECP256K1_SHA512_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp256k1_sha512;

localparam int TEST_VECTORS_SECP256K1_SHA512_NUM = 318;

ecdsa_vector_secp256k1_sha512 test_vectors_secp256k1_sha512 [] = '{
  '{1, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 256'h34d2f1a567d7e647b178552dec35875a2cc61df3ce8ae2c1357ea8c5ff505561},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{2, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 256'hcb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{3, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{93, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 272'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e90000, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=272b(34B), s=264b(33B)
  '{94, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 280'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe00000},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=280b(35B)
  '{98, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 272'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e90500, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=272b(34B), s=264b(33B)
  '{99, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 280'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe00500},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=280b(35B)
  '{114, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 0, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=0b(0B), s=264b(33B)
  '{115, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=0b(0B)
  '{118, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6eb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{119, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h02cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{120, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a169, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{121, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5eb60},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{122, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 248'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=248b(31B), s=264b(33B)
  '{123, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 248'hb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=248b(31B), s=264b(33B)
  '{124, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 256'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5eb},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{125, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hff6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{126, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 272'hff00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=272b(34B)
  '{129, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{130, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{131, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h016cb914246e1c92050a03d9b0b4f05dde199ab6bf23cec3a120f56da5843de32a, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{132, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hff6cb914246e1c92050a03d9b0b4f05de0a43cfcf1c53d8329a150b08be3d160a8, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{133, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h9346ebdb91e36dfaf5fc264f4b0fa220a11426278b79dc9a9edcf0e74bf85e17, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{134, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009346ebdb91e36dfaf5fc264f4b0fa21f5bc3030e3ac27cd65eaf4f741c2e9f58, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{135, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'hfe9346ebdb91e36dfaf5fc264f4b0fa221e6654940dc313c5edf0a925a7bc21cd6, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{136, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h016cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{137, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h009346ebdb91e36dfaf5fc264f4b0fa220a11426278b79dc9a9edcf0e74bf85e17, 264'h00cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{138, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h01cb2d0e5a982819b84e87aad213ca78a348979bd990065db64a261453a11c2d21},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{139, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 256'hcb2d0e5a982819b84e87aad213ca78a5d339e20c31751d3eca81573a00afaa9f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{140, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'hff34d2f1a567d7e647b178552dec35875b7217410d1f42428575ac4a392f1a1420},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{141, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'hfe34d2f1a567d7e647b178552dec35875cb76864266ff9a249b5d9ebac5ee3d2df},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{142, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 264'h01cb2d0e5a982819b84e87aad213ca78a48de8bef2e0bdbd7a8a53b5c6d0e5ebe0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{143, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6cb914246e1c92050a03d9b0b4f05ddf5eebd9d87486236561230f18b407a1e9, 256'h34d2f1a567d7e647b178552dec35875b7217410d1f42428575ac4a392f1a1420},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{144, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{148, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{149, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{150, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{151, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h00, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{154, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{158, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{159, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{160, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{161, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'h01, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{164, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{168, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{169, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{170, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{171, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 8'hff, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=8b(1B), s=264b(33B)
  '{174, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{175, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{176, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{177, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{178, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{179, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{180, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{181, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{184, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{185, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{186, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{187, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{188, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{189, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{190, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{191, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{194, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{195, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{196, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{197, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{198, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{199, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{200, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{201, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{204, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{205, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{206, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{207, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{208, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{209, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{210, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{211, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{214, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'h00},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{215, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{216, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 8'hff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=8b(1B)
  '{217, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{218, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{219, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{220, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{221, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{230, 1'b1, 512'h39480155ff8d0790d7d2e9ad2adf5513477af6cf22d1be2450d9b6c0d974c6a0e75acf16919577232616f6b835e80a82529bb2fe1065f2d8579e71f54a9c293e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00dd1b7d09a7bd8218961034a39a87fecf5314f00c4d25eb58a07ac85e85eab516, 256'h2c8a79b49cae4ec15d293575a5a1af5b4d6efb74ef5c2c1be34e33cdeb7113cc},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{231, 1'b1, 512'h0000000001b99889c891f2468c618149cb6865b933cca31eddb353de09746b540616ba69c5f5ff992c6d6177427daf1cb46a4c5c08625263a615fbf3eeaae178, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d743c5d76e1193a57438f1b43b1b0e33d0d1ab15bd3d57a5cf6aebb370d46ce0, 256'h7df27cb730b33dfe01e34a0067e548a98c56846d9a4cd64a930c96bfd917cf08},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{232, 1'b1, 512'h7800000000c52e48c315d5276f18d994c345b5805aa02872c29105d1bf75f152042a782853b4a3850822714434fefe3db00a19bc7eb84029869a7c1dca47ce71, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ba30f4ddf3348f26835e9c50f6a2d5023a9a1f5fe2e9cf14b3270015dac283fe, 256'h1d1616abb204f615fbe99860d89158c3264182d617ac9f1560fa8291b349d579},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{233, 1'b1, 512'had9a00000000987c9531c475b0236659fdd3dd795473bafb8f0753bcaa4bea4e6418f79cba317764c48fdfd9461986dcf668f250be9ed2b7b75afaac70ccf0ec, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h551d72e63f7b27283c4107f7d851f387b60f3f4713a5d35c21fa332fbeed4494, 264'h0080914cc37a3fe13a74db7fcc5226388d95034a50a89a9b2fe9bf42ea29e5714d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{234, 1'b1, 512'hb3284200000000930b8b98132341f68419e3262a7f2b8d60cfee7e1e364b36ed4f000bd5fcde187cde7397820b85a174025e4d54d70cbaa80d160fc9cc72d56d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0080cead3d165ce05c7cf8469f1c35c5a3a641696c843bef0f022a6c68133dc49e, 264'h00ea8409d743a4ad5e136207736c3ad79c8cfc7b57ebd1bd9b8a596670ad12d41c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{235, 1'b1, 512'h3bf2ef06000000009638300311c31a5caa29197ef0d079767e66e50824e8d41e5a36f593539a6c0ce102a92493c18061c70eefb94903831d9b8ed3291d1b9829, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00bbc0e8b7721065a51bac9c3aad64168998cc0efa23298340d436867cc86ba847, 264'h00ae3baa131a83153cb31de2f758e45139f62fe6cc9ce3941c6b1789dc1010f3e2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{236, 1'b1, 512'hef200f1a5400000000399e032faaf4b3c32d804555abf20471a3a18dc46f3917eb9072220b5d5f994d27b221346631c47eb579d69cc5e438b7e7b963bca9d84f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3a5ba93917b954617b40e1d866860d1522b0d310cac2457636e54e2ffdea888e, 256'h3eac6fe762aee127837c2c65fd9c1f65b404b2c31bb945e75d6166503fb5c8bd},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{237, 1'b1, 512'h7f12580858d000000000055d6877381f726e0a9237d1c012c9840b5b3fbeb6f43027bba37a94ba5fc0dbab436b88d4a7cde6aac151b06214a00cd8fe5f0bdef8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h647f2b4bef6d1ea7908ac5f3dfd705494c2587456557805fe64a703b2b17503c, 256'h20e164bbb505c6df56455908008cf9626df320f48aa3fc9d0cc8ad8bcf078cb2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{238, 1'b1, 512'h6b4185d1e7382000000000c86f684e5386df6f2e7e1dab4d1be30ccac1ea33d4e82d455b12857120cfb411b75c8df08758216dcb774dedf1438bd137f831b27d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h008aa653cfa001798c471eea3199dc975a4dea4f7c1ede47453409e606d05ceb51, 264'h00cab20967a056c0ea7fe9cdf8e1980f55b1597a2dad80c9223a0fab15c314fe6d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{239, 1'b1, 512'hd40c1a66696b7a6500000000ebb22b0b1f80b394770ad61c5c42ff0584ed4c84a3d185d3c07725f0d3080b451dad86945cc9b0801c01e0b6b8739ff8ec36df22, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00842e421f33be241d27f12f875355902a25819f210b3685ad536e23594012d9d0, 256'h4fb894ae0e9c24b6ed280e224ab0811469296a9837d1e95b5d9d661d21a1c255},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{240, 1'b1, 512'h68481d736990000f3d000000001bc2164f3bf7a43f3c7f23a875b84fcc1d1395c9bc3eec02e9aa7d38f4462d5734ca53f0db4e46498d1b8c9f9f4c92f4fc0532, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0b703fd75bdd8dce4820fe130a0b0af17aad4e4681b0254864d5d6f8931ff573, 256'h404521acf84e72ff22c2ee05d14a4bc7b70e69adc78caf81350e01379694c3e8},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{241, 1'b1, 512'hcf9bb31b573fa12e7e51000000004b37d8761e5d50f214b30bc2b134bc7e0e30653b8debc737a21392357313d13e08eecfdefd8d37bec92b680a84f5430fb57c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h62f0df1650560a5800fa670377a4317a604d6475c490066ce15638f8d1330b63, 264'h00963edf905197096818368a993fbffe32908a57153e6a1612bae6ee9ee8a8a719},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{242, 1'b1, 512'ha678a93e12f88e59d6307e00000000bcef462484d98a07578e5106f6b5e6cd1618aa82e3797b4bf519cdc4704616039255cb3f05fc8b93e4a48e2c4cd5333450, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2901ade694d4b9c376b3244018e57bcde7057e8e11dd0f7d07080cdd1a39194b, 264'h00ee65a4c2baa70f8e236ceba9eed400d899f75276f94e4b7997b2b01ac008bbbc},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{243, 1'b1, 512'haed2cc5334773206d7170bca0000000081dafcdf0acf2107d7c016b54b1c0ef3663c5ba78277a328ae547ffdf6ef2e385a374d9355022f24dd05ff9b357e5039, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00aa9c8e5311b232b4ce9db03892f26eb77d655c6ff09a599424abbd4b11e750be, 264'h00c1034c44b02e2fdf05e1ba5eebdf954c5a01794600059e05e5c73d542da3ee38},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{244, 1'b1, 512'hfeac570e6cd1481ff79f34cccc00000000eb127fae412cf598abaa6550b4f5f2e1537dd5c5d6c57b0b52c103ec0340c9e292d0a263d74e44301efe65d505ff9d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2febea016e55059e91e157b988f86048db57c37fd122f5cc60169ff4fcb4863c, 264'h00eb19cbc35b3061e1ac4b59b92d1f732cea3212dcbe943ccad82d32740bc22c33},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{245, 1'b1, 512'hbacfc820b1f513e6a157534762b6000000008ba56a4c814c4c12a828e658c8f7d0453900871cece52dca13f4f1df23685d1bd43488e2acdda903b2e0f72b9d64, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2be463ff06af2096dd62f0326e1af51c585f18ca8f8aa361dedcf55d543e6b7d, 264'h00f56afd59dad42530d94f11c59a6408c54826b7a9ef83f4d020f209d71f9b74c5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{246, 1'b1, 512'hf9f58ffc6e2662f4992e06774f928d0000000084b7ca7f7b6fb750919f466be3366746484849f67645a424ce6009fc560031052d0775f47984d3a4727776b916, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f61f64defc45abe284b39161b49585f21edef1e88d06389e5b5aacbb394ce4dc, 264'h00a5a27e17df10aedace97eb2c48659f69b58cfe76a1f1ac30fea3043655bde515},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{247, 1'b1, 512'h5f6f67fd931001c593ff6f8e5ea8faac00000000ecb4ce9ec81a128cb55bba07a9b186b28f7e787f7bfb7ea32d9047b830a99f2ac4144ee3f6e07ddf00e68646, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h052134eae13c1dec5ac5aa46186391786f5b60591cb0dd30bfc61e89486abfe2, 256'h09cdaa279c4f0d3d5ae00e0d74e733a260b8b120a1bda7e5a90194ec442e592d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{248, 1'b1, 512'hdcc948cfcd6f3cd3760d678a643ab0ff010000000095bdd5dd5c0b9579c7c6b0f3e921033117737e31acf8ab117b62ee54a25abdba306c71bb0c3d60097a332c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h24824614686b80f3b738970a27816f58cf103c4a93c2d6b0f5f6de65a65501e3, 256'h180e5801a593063e75b83cd7ab8e52575a013a1be5cdeeb05b30e3ac9dc4ed82},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{249, 1'b1, 512'hdfc50d9e551fd99c3ceeeadef83e2fab3f96000000003206a5e2b462805d83d6ef6280540f3bfbb229421d6f5f2794f117259f9dace4f82dd57889a74a0fcce9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2ff7a5ab2f1a3323651a0d17c4263672ee4d2c560cda94e7d52ee755138bb045, 256'h542ce83d8d9d441357e24b618b5695164d4391791cff62eeb01609d1d7cb1c0a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{250, 1'b1, 512'he4edde495afeff435a69e94a6493e4ec2c0b1b000000004c8e512f917698225b0189f732d3deb6d8c1c39b6b59e0701bd7f7605a521891358603454d151d8e7d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ae446d1a81766d21dd7fc515d0a956605d0cde26d6086a76f8ffc81a6dfbea46, 256'h4fccef9f75e94abc7eb3f2bdcafdc5d97d61b9d950a06010ab4c54e3da7fd4e0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{251, 1'b1, 512'hdf8f102f7c54ce2cb6ca609ce724818f7621cdc600000000c69bb15b7c33f6b27c75a153b581d47b99de18ccc8105fc3bb697f180112706c5ebfd6fc6c8a6322, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3957cff4a75fc6039c0b0c2e47eb9b07ff6ec5dc8a3c3316590a7ec9a1d7d993, 256'h4e578ee6594a00cb80c640cb9589d616dbd1cecda2d15dcc0062f30686d6073b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{252, 1'b1, 512'h3e526c3c1f02aa2e007cecd9e02f7dc3d06f361a0c00000000f8e183a89a7218d8183a928d91c6bba47d950bf841396e5fedf9d87f66671deb8d2ebf63e39751, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h437c36031737a3140dc30eed281adac8e9074187aad41502a3b9a3bfd4ef252c, 264'h00da13f88f633202b9b9517b93a6c08a7b8e6858734e8894b1a64c6ec08f1d0423},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{253, 1'b1, 512'h7a750c1372a8d9b00991182aa031522b94a1a7f4509a00000000baafee68e65ef0a94f7983cfeb9241e0b7d8fd590a0d55b16041eaaabc38e982aaaaf6eb75e6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00828c12fd9fe31f91bd8f58aac72ee6485e34ceddf91927cf3a09b63363b9d8e9, 256'h0e889664a8c98619cab572687064edb4f0500f8324a5df0bfb5a431a3cb1ca39},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{254, 1'b1, 512'hb8df763eea0cf11e9945dc5667b0147cf8684d618abe1200000000917eeb543a4dddd7217ba71e998bb9c5fd62b57509b7cdb489bc3b64f66a70e4b5c12ffd2e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00807cb34aa6ea48b175f41f3afdf70a109d2b746ae48e08677cdafc33d916b2da, 256'h41980e6f7ad19944d278851f98e0a6220ae888964ae81a667a63fec21449334d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{255, 1'b1, 512'h88670299bf6b255d331cd40c7154c438fab9fdd2b4319e440000000057a51b1cdea2812fd594a8cdd56b4f5cb069625524bd53a5f304653824d4afbf9bc58d02, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00a998f9f0daf02f717f5292142dca447c722d2394dae0c84910433754669716ac, 264'h00826fc37269539cf8a98997f8a0268bfffe888d6c23bc68ad7c759db47f65a925},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{256, 1'b1, 512'h295422dc27dfac13c79d2028d3daed64c1dcaad525dbbf14a9000000003667b1baf41fd9137fa0bd8c3851590b206aefb6cde62fb4ecc23ae308e540e83a7f09, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f151b614afe5bc9d511d0c34a7eb44283921272e91b3e5d02821cf7a43a92bc5, 256'h097aa33dc50ebf8fea036cd7e224a4d38aa20773e5a78ddb83a2f3b579b2ef6c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{257, 1'b1, 512'h118422376e38638a08705cddcdd319e26fc8a2e6d4a4d1400fb70000000005687b339ec07f51592f6e254c9b7291fa2d0302df9fb2702857e3f69bd4fba01654, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5f21585381f5f42e9f76be3f61f4cfd6476ecc6f06cd4fbcf13e08c27f426148, 264'h0095d5b2deabf19891edd41ac52d9072fadebb2f0145bec9b916f68fd1fbcfb3cf},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{258, 1'b1, 512'h5a4801a1f7ef2afbf8e0e76cbd6e07212568cb47638e22e55f8e6c000000003a2aff81ce04258211030942fca855cbc0ef482027b17a7ee523b15483afd91355, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00bdc361e68984482d7b169bc5e6ccf82d2263871be749d67a44f548d32bcaf5f1, 256'h375614fa4134d5055ac117a6ea948b74269b8063e39259d494a7544afb6291ab},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{259, 1'b1, 512'h057d7524efbce651b92e0a70e4454156e7cd4b696c197c6a064032c100000000768565d4af2019fe3247dba91948292af777f107fdc9c3b47659eaeab26ead77, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5773b016dffac865ab008abe8a06353d197b4dff32403d7ce98ada4d20ea8a00, 264'h00d60de9c98cf50eff0515b962dffd6aac8a1b72bc9cfaf6bda12b99f63eb976d2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{260, 1'b1, 512'h31ccd924b687a2a6b70f4888ea911ea38a686e56e5540ea692ca3174bb00000000246ac69c46506bd8fe924eec33b33ebc9f508d4251c459fdcee3b4c84d4ea3, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h57b747d21fc898472a888b88693a989eabaf143396e4cb2de4af19386fba384f, 256'h7c99f63904191a4464d0d23ca560d5558895cdcff93af4b00c1c66ca2d974393},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{261, 1'b1, 512'hc7b70cc4a55d55342487a4469ad2243ef6d6b69f11604b8c12baa03dd3e10000000014df0db29a9d4d54b26f4047f3e0c739f7a260768b20589254e1235fc590, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00854be2bf302a2d6db437eb9e78703673c1c7371399e68caa8625bb13c7aa0fec, 264'h008fd22607e0169eb2e2e00c4af898fd2a609dc57a9fa94a7f93372098fa675649},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{262, 1'b1, 512'h1634df8a3271a99f360e3bbdcf789d24bf4bb03e3114ee9f0fa930541f1ae0000000008d976fb74f27eb316ce3a24d92a53833e600c353300f5c4fec6b28c581, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ebb3359de3b13a518545a86b7fdd92f4793225b8ca4555a6bd4182922b0452be, 264'h0083faa7dff1aa0eed89a7ddcdaa5d716ba6253c5c21f7122c2755eb78b28884c4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{263, 1'b1, 512'h8f90b6a8ecbb870dc24832b1f4719aae2d8eedd7faf97848b08d2b528abf5f44000000008877a6157344e6a9dc43b90c8e2dd7ab9bdc5237c912e094660d0878, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h008bc91cfcfc85ba8aa171b703a330e398df4460d22602e73e327423ebf98bf632, 264'h00ec7569072aa73ff19f183daf433abff142d7d5edceb25b771d853acf0fbd68b6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{264, 1'b1, 512'hc0891fc626ef4b106fc00f5c067253f26a2868d09aa2ce029466f353ba525e757100000000a3cee37421995445fae741697659a406394c870d8bdda130080d15, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00895b07c0450ed6f4941633a053c978128c46e5225c00eb009c3c6cee5eb2b842, 264'h00c982818b260f1650e03eba8f9db1a2ca79c3f804dbe7d172233260e1a9c10640},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{265, 1'b1, 512'h76527097fb3945436a30cca60392c170abb7ddf6ddae93e3ff7651d468eb3e14865700000000bd314c31706f8e4d1d853b151f5afe680e13cf2f255b2bb697bb, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d5e152ec304090d764fd7ae61abeeadff2fee8df3dccd8fb44d2af5a8dbee0bc, 256'h72518dc1ecc993faadffc3426594fe2024c7c84ba101a9274d88009393103ff6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{266, 1'b1, 512'h41d43cb27d4db522756dd682826eee8d0f60163c7f3ce67a39d89d7d89e24818c354ef00000000cab56830cd18f7bb9a7d1b2440fde06ce647518fada2dc988a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1298b131ce97a528e5dae05d92b286e2447b17ec002267b9e8f03784d4074bd1, 264'h00edf223ad9c308aef22e1e0c24a20268f966cc2b9ca4d941945bbca057db92d4c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{267, 1'b1, 512'hd34ac40ed5ab79a4e5ac1e4081e0e47e4fdedac1555b01ab62a13ac0ae9dbc3c23f799510000000010116f328ad1db0cd68cd1db9e1b34b5a52ebe9b8e372b78, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1e79b3921d23d290a57d08958d3ad8305ec444efe1281c98fda44e8af7648f49, 264'h00f4c7610ad1ba9339178c50e7979b5aa9af07d8143e59d13a2e84f98f37101e3b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{268, 1'b1, 512'h8b5db6db13b1f5e609965dc38215d14ccddf66a9d86505a67cca37f13cc420803c1df80f4700000000b044bda09a83e4331aaff90c4faceea315e467f5fd91d4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e455f464e0edff9c959f84f081828896149a330361ff2d16d5a2448c9d683684, 256'h351cfa2f29a1318ebb3a46f0a36df8954043949b8d7cea94eacf99108b4d3fa0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{269, 1'b1, 512'hc771e022bc376ffbe1f513bcff11884e790e53878c197014931f6360c517ce8de1c059d091cf000000003c560cc443a6f005ea58917a52ca9bf60163afb16ce8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00a885770c9ffef33f0c11245064936e3dd165ea2633575a6a155368670351f726, 264'h00de31e6a58626a41fd029cf766ef44b8273b88558e2452e893978fbdda1e321d1},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{270, 1'b1, 512'hd9cb55a3f1ec161bf6caf0452bd6d6c876b35dd1000eefe18378afaef6280348fd799e624e573a00000000085b3b24635f5c10770090ea935f198728655e236d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4b6b451478ba253ae3c75ca5b18b70ccd3cca408ed245cb2af3369548dd2e507, 264'h00fe479b631a3431b42772925cbfe8e789f9c55fb2fd1d7ab51664cc2fa571ad93},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{271, 1'b1, 512'h0caacc1f43ee27ec7ad5269155a66172ac310d4e202a9b7d3defcfb07ea8da85415ac2b116e665830000000009887d6c7da6cda824528345e14a6675de23988a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7ca70376547ad6d18f8e539f09dc269ebaa06854c1adacd58fdc735ed3cf0c16, 264'h00f47654f4c0ac1b0e65b712300e3bb472983b116db5206520eabd886dc706b266},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{272, 1'b1, 512'h5d761de2a231df86c0fdd90da20e5811f7bd9bebb3f1966359b8fdf554f79f0bdd32ca06410e70e61100000000ed3d4140a60908e85f7fcbd26dc792bedacbfa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h388514d147664fbb37271cb8693e47459c0627d6b1dd52dff1d3947dfc9cabec, 264'h0099d3d40814aa177be99e4819696996bc75073f4518955587cd56b5ad8bbc2c58},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{273, 1'b1, 512'h78adfad2734b7baf32f4e0201bd6c3e9f6c1763cbe35858a0f56466db34dd98a0fbf5b2a71afbcdeebd400000000d3da1a5035406b39aa13c126a3946b6c6a5e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h44d3ac50d9b65601d79b47d6c5d98394cef155211ff37d4bac15e0d4890809b8, 256'h3ea03829afb0545e088361a8cf952aec17bab7637fddd6db35f039803523c921},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{274, 1'b1, 512'hf1d6ef224f72b83a109944afbfb34ae1f70d6e50eee54a91faf8ba0fc062563113d988f2b826c055ecc61e00000000554878a7e761e75fdf1ed2ad2d138b2974, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00a33004a2cd50a4f70447fd382e7fdc9257c4d9be7b16e686c5082a231ee7b010, 264'h00d87b96ed3beea54652607017702cfce5d4e7fcec1fdd28f41681ab80a5c5b63c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{275, 1'b1, 512'hb33f308c5b107050cb2e513fabf8b896e52c85852fbe32308bee8b8661121bdac78f52f924cf3d5690ac92d5000000004f0f619e72ec1464166078ba3f508a66, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h668ad18cc22c1d1498cc8e5a11e2bfc4c1e1fcf0a7350a5806c5533ae332f0b1, 264'h00f58b49369771bd20bb08b63d4a9212e2dc71da9257ed3710d9eaef9bee469eb2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{276, 1'b1, 512'h0392f8c2dc961605c5693d9452731b6a8292ff57d6995aeca0dad3117459668ec7809dc09cf154170fcd624be50000000026e3d92dfdf1a2abd09392468117c9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f7cdcb0281c70786cc3653820d1756a78395a9eeeab2a4d164e260f64ebfd6a8, 264'h00d966c74499cac97ca8ee67400df01b14793b6d7d07668fc202a9918f3c046e9b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{277, 1'b1, 512'h9dda0539bfe47c75bc00b014dc6046c9db5d7a5723acddaccaf2aac7a9250b732a80cd948409f132d1dd65cfe91600000000d53c76be9f75fc6927f818acdaf7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00de0e781d9e3e7f73021458fc1201fc021e5c54f1fe40b1b10db8fcf16ef7e54a, 256'h7d9db92321b5e5bb105990145390979390d32394116f4e78af34b85105dee8e9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{278, 1'b1, 512'h572e1d736d78c42eed5ffabdfb25b5c7908aa60728ddb3d36a24c285db9ab996433827aca9e23716c3baabbbb4527600000000b9c1a728fdb6f65c10935e9514, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h011dac8ea37f7bc6a530a42d0e3bec8c845694f73bec6950081a6f999ccdfbc6, 256'h153e57ee45e0a379839f3b8f6faf86de7a626b210f4c1007e431f842e39bf7d5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{279, 1'b1, 512'h81b675425e8c528a0a51b23413c8b796411a01b207e0bafc5bd2a46b05237be84abdae1ebd492fca053bf7e3133392720000000086ce63108f1dc5a3b34c575d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h63f9c43a8cab49f518685a120bd73a4e5956f9f167a78d4661fc795d41be2ae1, 256'h6aaf4f3384f1489ef026cb29e97ea1b5562fe8ceb9978d506fb7064f427b9f31},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{280, 1'b1, 512'h11c203ef3c8978266a73147233f7c9c9d16108a07847ff587f1e865f28519e7a161664edb56d9e791fba0717124717b3c90000000013c59e26ab63c4a99b871c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7f0fd3736166195ba810d5a2dfb5e1f03aece2170510c8aa4cc4a0c974a7c5d6, 256'h370c8772a75d32e8c9cc103004e75e6d30a8ac8611b84b89c41c65542171bc5b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{281, 1'b1, 512'h5de83c97136ff31a90ea5053ff256d522819626ae3734c460ea7681fbd0a94538ed840f3bfbf8055756e761d8149786b8cb000000000f37f36e4d32d46cb9bd1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f975196086d10f683f4aa1a3c2d5fe13fd0f52ee72aa3f785006aa024c758735, 256'h6a66364156ef21b5dfdcee60cce8fb09c12019bc576848ff73db49856af74681},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{282, 1'b1, 512'h4a5e1e8c073ecb2832fe0d0df42a72ce225ea97ce093ed320aaba00cab25ec3e90a6aefaae72ad40273d7309e40582f40a37c1000000000b1e8576da0eda555b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h35fe6d9bf9f7d47612c3f5be6a4e9a0fb0c14854d1a377adfb5485d6e3835c6f, 264'h00f96587fc460e7d07396f9f2d060693dae632721259e77c90b8314002a5235dd0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{283, 1'b1, 512'h9f920bb92b4527d54ff6877b80c81585dc4d3d1e96fce780b030f9f371f8a1b68e2e7a86536acc3ce96737bd5fba0ff669f6b1600000000000b5868a36cfe6c5, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h210c7c9b231293c8ec09b0f610d31724a045f6a33f84423fdd541ac11ff78962, 264'h00e5a40e6b80da99cfc49ce969f1f59146835183e61001b4513f927b71ec3b2a13},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{284, 1'b1, 512'h99f941e73ab790b224ce0a799133f6b04eb9bcfb2fd0ec84b8e7d5dca6ca50d2b1ae4d31c57e2e54f97f59b6a10d0758cfb3e46500000000909d4fabd9d1962a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h09b7dcfad2c84b89825cf3aaaffed51664faccc0d171a43387a6ff98aa128a04, 256'h272b00e6e0917afe4fbe782604428e09fd91c38125d51c3ba06ce3198e6bf736},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{285, 1'b1, 512'h202e258cee0bca789ccd4c29f3835362b6f1f53faded0f1d58f4ff768f6202a6de3ee3b922546127fecfdf1c0446605751df9b7fbb000000001a8a11a3e383f3, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h09c7c99681c9159b22c0a467999559a31e279075d37ef872a88ae13565f6149b, 264'h00b0ff953be1940d2cf548663c1b4db7b416521db289467733b9a76629f8ab261f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{286, 1'b1, 512'h8c4a184638926ecd8f6ae279181f9171181295757e3eae5b5a0de2fc0281358973a355e4820da4ce0c69db549c72ea007f80ae990565000000009e51983c039c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2bfaae0ea6d8baab3e02ad7fa3dda3ce0725d11533e3666477f54d697e2ca9bc, 264'h009289d5da443395bca18fe9d1a4afbe04a32b4ecd258eca6c1772acff2d0b9a89},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{287, 1'b1, 512'h92eabef5ab4296dba863345a2f11c2bc8d32bc02731323a19a88897aa1421f384448516975b6397a8e627fd3cb5a5dd6ee3c50226b18860000000077b18d5c83, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h368846edc677ae8fc237069cda719af3d7f17cc136fe443b2af614ccfb4844ab, 256'h5ebe6c1d3e88bc4e291841ea97c836bdcf67d9eabe926346c5f42105f7b38f67},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{288, 1'b1, 512'h4cb05f07197bd719557dcfbe1edff395550b275100cb073ecb4a0987621f83a5f041996f63fececb77a30cccc5f8067e36f650f7defb611b000000006a949e2d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f336da82bea2a111bddef6a25de4ab87d7c95aa80d21838f3a4efa3d9346555d, 264'h00da5ab612b327aa0fe95d1caf85f3b6698c23a47212006c5667cfa92aa3ef4dad},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{289, 1'b1, 512'he744eaf4e9c4c17549ca3907721df98de95b69d07d56eef509d4740a3cb142bc61b6c4d108676526d5a77188977d924dc9a8adf6c01adc35d6000000007f3077, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h0097c2fb9865f9e76f8d54ce957120b68ccb04cd3183dae7130f73139cd56655cf, 264'h00fb63e38176ffac37d0ec1e49c2e2efeff04dffdad5a75f3576f8276cccee9851},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{290, 1'b1, 512'h4fbf285c9be6083627ef151df0d2c5fb00b6edcfc44216a30467a4fe268214ab66dd9be898bea57b48f6499d09d4beddb7c9e8bd813fe7c1cacb0000000054f2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7393e0207e07bd73b674d3667dfbc9c30022574d63079a040a23c0cd7e1b6aa6, 256'h2994b3468432fecd0a32134171179d2809244d586bd971129cdba73fd3dc8876},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{291, 1'b1, 512'he698cebca57a541614e179f28ba51cf82fa0fb4300f81df5fe22b635eb4441b496a36ad280999f503edded3ae1cab1700758b5ae80ce33dbf25c7300000000e9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h21e1943d7d396a8c46658bede4ce155c9a06f929cf6ad292d32c91cf8f493887, 256'h30783c682cebfffec5787d762bd725bafc9c4075ad8eb1582188f4c05dd5169d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{292, 1'b1, 512'h43f5ecee4c9b5bcf2497d9753beb1eca8a01c143f8b50518e83bc7f3f62d049b03430a6dbc9236d54b7ef5475a232e3de9160e9649e3c8f46d2f1f7900000000, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5a269eb44e910bfe8a2656dee47556cb908a417917e2068e20d201721f44f9b1, 264'h00e69d463204dce77c249439f22f77cc4c88134012a286b36a9559f694203766c6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{293, 1'b1, 512'hffffffff4fbe152fff953f198736b155220dfe633b6fc7aa5bb392cb96cde9fc658b17828d0d04ece0f6e35ed6bbf357b86665cac7735a3b9c85c038d4a85019, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00cb8c146fb3d58846e5748c48742af2f1b77805f6cd1e4eb98d8c66cbdf5d6455, 256'h17ac992e10251e334467f8e57e2e1c269db8b19469321c74b443972a80f38b2d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{294, 1'b1, 512'h47ffffffffa19c2322e79638701c393ec0df74b5d27fb9ea7cc3e3dc8badffcac83dd8c409a22c2d7a64b5693f153f60264487aabe5df546115cf2eaae415ac0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h212d84a153db81cea5212fa7dee31d59bdca1307277a01b5936c3aead31bf1e4, 256'h520305dbef2bda6526fa2cfca789a1c9aca5c2ad4c0027cc8cf3881813da8a72},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{295, 1'b1, 512'h391dffffffff5a981c0576acae266e7b35ecdfeddfeb6db903e9f4eab200dba039b146517f0c5b418d096addeab6d0962a6f77c2a2a552748b788c07796553e5, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h310c82892f571134a36725f4a31c5cba8bc46e65002d73b11364084433d8da4a, 264'h009ca552aca84b96cc9461e2b65a64975118ea78b8b355a0ebcc1a61de37877d13},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{296, 1'b1, 512'h8c8ed3ffffffffd5bc0cf4859c831b89860c28ba17ff5a259b6982325be66498c4ac3119da331db0976678878c73473aec528a7107d0d9b1a17dacb9a9237b1f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h489deda580c62533783df9fe62de34c2e2cab91d676709beeff13afac8e90db9, 256'h32a85a9c56f308b7a794dcce614a5ed7e0857030b8429fe3b4e07ad533a5a00a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{297, 1'b1, 512'h531341a3ffffffff263c81971e877fd7cd8308b0d536d7fa3c88e3beaad332ef664f76387e4c43dee6c0a06423b18d1b1772f65acb4f9b672b97a648cdd25929, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e8897c1cad1fc870a7d364676a9d7f7cd3ac951f3bc3a9ef1f7231466c3493d7, 264'h00dd2128e876d62da82cfc5fc508d33bf66b71c0a84d0a9b7e47dfc620f5846bc6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{298, 1'b1, 512'h2639a8ec01ffffffffb54d98af88ba2ae383d69bee2f5fadda599d58796fc766130e3fb8f4ec1afceb8a1c1faa3ad305a0fdd65796adf8ac579c1306d5f0195d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b4d771d19fffb1fe5ead25ef5dbf6b53d4d3dad284641108ad84b2541ad435a4, 264'h00843ecdc2641b33a3ae9ae15d559f6229d7304ee5ecabe00db73bf2b6b5c6c21f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{299, 1'b1, 512'hd9753a5a8b1dffffffffcac9aa24c9d687a2088ed837789e72d457d0bc67f54860087c3f0509744e0b461f88893e2de6c757705670006c9e9e8c4c3757fcb160, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5ab5fb3136fabdbd22009642df03685935819895d675fc284e8b8112db522d08, 264'h00d87ec88173e823ed70438fb1088b00689352542fabad5e9fd6d4c3c58f722f86},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{300, 1'b1, 512'h9a6bf9edc61a22ffffffff703f4706318ef947658ec44c90cc1630c916924f1635efd88bcb900db41dad160ea33f8176397bb8593e19199207ca7d57bbd28305, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00be310120169f8d488c6e5ec5b5e588ab8a65040169d9efd3062e0d05fd7d58df, 256'h45033f291fa21a85cc08f78fec2dbd94135520de261360728b8743b558ed16f8},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{301, 1'b1, 512'h4c18a4947b15af08ffffffffb9de1de3873b4c26280b1286a51715dcfd1242208ad49b2aad0864d5a4529e4a653d7a6355b7c1747fa9d876159d43806661395e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00cd7fb3f2c25dfab6f9ee83fcbb08698680e9d1f3d47815bc772d717a764f9997, 256'h287dd85b976d7f56d23ae7837398c118932aadc982f675f94103036729a47c7c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{302, 1'b1, 512'h6e50953fea8dfead2fffffffff824e02147d010595358c98ec376055cb9ddc1dfe6d3874cf38e8a98ef0664fd3b10605bc14506eb7e46460c9db81b10e2f6730, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h69f18c064ad2683cc1b6d8b79020aacd186b6ad1999e6e55bf28bb1dac33f339, 264'h00ef66e66001fcc219c9a927d7f0b84863483bfd1ffa6086c06921905310c793e1},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{303, 1'b1, 512'h1539fd34220ed16ae0b8ffffffff88a04bebde47a3a94f1b86bc687c2ce7648caa7d42ac8693b5704e401b7c9f4864bbafe3bcf761d862739eaee02516a0d707, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 248'h547c6bb40f52d207fff796a29f6dbe62058e50fb73bde6b9c6ca11346fd8e8, 256'h2bc82bd3efc9febe8578acdbc3148bb46c41a39be9ae1994ad52d8bf13195d09},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=248b(31B), s=256b(32B)
  '{304, 1'b1, 512'h69e3c78c7125bdee7184d6ffffffff274929ae7dcfc4692b84880a518de1790a758005ef7d4e29377cd891eb08e9fda55ac99a11b4dc9a15ceaf8887ae941fd7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00a80496adce42e7971ebe91300710cf4f535fad266668d76d72c95fffe4d42570, 256'h0d4338ca32857e14e0ea8026bc194227b910b98509c8c9307b0d8d93d47b191b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{305, 1'b1, 512'hc3b630a45b21b937bf78ef4affffffffad33da42317364a1090ed4446da7738caefc807ed99c92f85a6f6ba946f99284d4b9793896bc5e0b6f93cf1b09b35a6d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3de40634d11a7a6b67023b84650420673ce6dbadb1159768cc0fd55f3784ec88, 264'h00a455fb08e51b8493177d88fca43aeff306e1490d7f6d24d6a910970a3d8619de},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{306, 1'b1, 512'h14f3b0fc1795c9d400d904ea0affffffffeabaaa40c2f532e33f6c61620d23188712a838f9bd1502b2a5c321117ed6007ccb48b375c581fadf340b0d7edcac93, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c1f229c0557d4c47962593781bc96cf745f3bd629ad85434dc2eee456ddb3031, 264'h008638f6c01c15d23db24bb851f6c63c763c1f040976f3f2b32c4bb1b9506c1c12},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{307, 1'b1, 512'h386b3f08bc91c7e18354f3d46de4ffffffffbf492f2bf174abad52337a99f29dda6891d96f85efb667480bcad7d2482ef7f32a314b4dd39576ef560bf01fefa0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h35dd4957b352e8b1bbc80d1deb21f9b0989188ade3fbe46f75106da1684e1d6d, 264'h008b508e2ed7a51efea0dfaf377f6bd5d4ae133cc4c93650600be545af5d3acd75},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{308, 1'b1, 512'hcd86d593a60faa34608d5bcdb2e878fffffffff06003c116f812eecd35fc6f3cccc1dee24c5cb89cfe9d41b0defa4e5d16b1d9aa4897e6efc838a8a6dd5f22aa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h410aa9c943e663082c6f76b84469c9845e0d439ba7ffc7cac0418eea0e20e638, 264'h00c873ab5c21c9f0ce0bf78484028796b77451e1187250ee33535dacfb3cee5f61},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{309, 1'b1, 512'h7939a3e06bee091634b535adc98afd56ffffffffeb0206c5b2cf892d2c8fbb5a2e105567cdc4447b476525488611a085b870e498a13b891cfb9a66ad725273af, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h008191db069b571cd40f2676348433430d3a65155c233c46a42a4299e6f5be806c, 264'h00f3679ef8af0b1b3a3aeaa7bcee51ce960441622e9ff2dcb22a8ec8de724e0a0c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{310, 1'b1, 512'h180c134c29d50916f2c3b32bf43382eeb0ffffffff6178b5edf0856813b75ccbb537c57758d3e55c190bd8e648a79c5bc6a62e45f2f037aeace1733bb7260707, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00889c44edbf3825b18d933aecd5ef70d12ebb00bf79550451205fd6f5ba7f372b, 264'h00ecb67194bed2b8176077622d58c9ab4fe4ca34601decc09f9386b8c4445c7224},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{311, 1'b1, 512'hf2694ba9c9a0d83faff7ff2f06f0495682e8ffffffff1d5cf19e626efbbb1425dd286e93044edf262236a46a82638145b4d15c18aa6e1edc919e22bff3a9c5aa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00aa87113aff2e1ad6461191241f90a23b91242d0066779daaa9506a4188abc427, 256'h33dbaac5ac443fb4d9529f83247f94c0ad1360d4d0ba8e162a377946c6ab9ae2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{312, 1'b1, 512'haa2db4394e6e52a9f0485ea08186ed648a109affffffff19fae34ae6524a6abf956c07617b15896bd3dff11cdaed4f9a2769cb4dad0b0e007b66c06fda3f256b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0e13f66a8ffd0da1c4b67f4d805941e90f98ce386540c48019c1ac1054075683, 256'h0cb489e8d5acfca5245d9292f59c6ede52425157af77b8beef38d23b6e6ade13},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{313, 1'b1, 512'h59ce78a87d80e90e1e6b70def3179e12e78cd5f0ffffffff11eee1f43a7030f096c301beb60d1fc2be04d27aaec7c385fb9aadcd6fa37cbea40783569080dffd, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6c1813f660c78bda956c1685bc924f69d1bbac5fadf3e4b027ab049bc82ad134, 256'h20de89ee005d7646f070bdac794ccce24d661b390a78851d35fe6fb5b25b3eba},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{314, 1'b1, 512'h5d07345f237708f45b49a7286977f331a27c8cc58bffffffff492a29a714f16596215046376e8d35cebaaa06b73f14ec0731a0607ab89c4edee5ad7f575c93af, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h48dc830b6326ec218144391b658d52045ef86ef918a8d41c59131912b1a46fb1, 264'h00a431916cb7cf79129b90f09842b3f2164a6cf603db88f2d99944142c00b42559},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{315, 1'b1, 512'ha6d55690f7fe8dc6a67ac00e5f136dab1f6855b53643ffffffff2585eedbf8e7c3db326f7fed8c48851376d7b1a34dfd79aa6837d19b05becbe8b8d122d1baf7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4d45782be145a27ae9ecb6cac1b9e30be87c0d13b7d6ada9f795ff051351ac70, 264'h00cf71d1eb15e88446ddb900f20d1e0739da499de9963fe99ded00a62da6462d62},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{316, 1'b1, 512'hd42f5eb7f42a9dd25a5d9513de8b6ccd5bbbd029263799ffffffff3baff5bcc111d8fb4f14fc4aac37a1dc5633df840644aeb69aa87f390c090e6730bade402c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h11acd8b8d736e7f00476495803fbd20ad351321e800cfbddbd6a7dd610c5ab8c, 256'h734027aabcca9487773dc3ab069b802c00f5b6e5520e7761496ac1e7c78ced91},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{317, 1'b1, 512'hbf0fafaf135ee4e03b991ef87e6e9377150ae255e043de57ffffffff10002deb92f4bf4c1770933d3137b0165ebcf81c8c3387c21457e0fe0c39c7c7947837b9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h41be8b3bf41a4c507de12f098f7d409a1f941fef84d93794c497f7242a7c382c, 264'h0081f7e7243116f24b84b0321e93eed35e2bdc32b00aa8eb9583be3e9b7a09a4f3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{318, 1'b1, 512'he0dff3b5ebca4c971f1da5a6726d24519e4ca71f45a548d85fffffffff415d9ea4bcfbe4749c275d6594e8ca8b76166fc90eaf2d9f466b0f0a5ed8c14eef030b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ea032ff41b061e93e456a5f0a9cdef36c0732df4d55ab4d3867484b0fc49d9eb, 264'h00ab298dd811826a6a9319c3632a96253c31c14f75baef536a645420442bab4d43},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{319, 1'b1, 512'hd9a9dae1785ef8a49d7c81b0637471693412a29484ea1cc780d5ffffffffb70ab50279ba56f6576dd87ea0cc08ed51afd395238936b4aef7284700c8d5aa9f05, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h008b1ff140c65adca22e5596ffb95a5121c356d2d4055f14606445249a5725686f, 264'h00ef8c16ff228114a7e33b35ad465f957577dea405fbdf3faf077a878754e58bef},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{320, 1'b1, 512'h75c7b98cfddf04426dda027ad897cd5ba9d5318c27288ec0f6fb67ffffffffb744ccbcda470681f3689c70425ce514d035e05dd133da5c2a104980f4ffb91014, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3a40e8dc3ebe9e19dcd0d4d1b698ab2a4934a146def5427b3a6a8fbfbf347846, 256'h54f65e36088d2d4543011c94b1e5371697202d488b342dd6f77a69944128223d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{321, 1'b1, 512'hccfcfe85e6d12e377ff1bec515ce149719d86cf3591b3dd8d4344022ffffffff60380790c2be6a944f31e63ee7b421a42ec5ab43f84f05aadc5ae5c42a6455b9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h15fecd439137df74820727f71218405cbe525d403c574471d8a36fa4b1f592ab, 256'h18ec290971ed0a227ec47f1e2142f3b8fe5b17336350c5515d4a87eb3382fcb6},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{322, 1'b1, 512'hc445da85686a33c8af5997da14f197df87bc3ff9f277b46831c87f8147ffffffff0970446a79a2c801e1a6f9c03509ae9b782a31b3b15dec03f5789a8345e14a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e676e84a299f481a207cde6a4271c87d73e29d1e49216393292323bcdc238844, 264'h00b8a98c769bf81429644758c8f803ddbedf81634e53099c43ad0ca42f4207ba16},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{323, 1'b1, 512'h6a94c0cd0809f1ee1c23039f735f24a0a006a0504c295289507a9dc93e34ffffffffd7127f6a21cd1ec975e05b1a8d78144da6293f4440723e7d6062dae06a1b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5116f8f0af12b47bd025aa6eaec5007d4e3c5a3a72cb4c331f569581adb01bfb, 256'h6962251da7ba9ac951cfbd2051bcb7d953005cb9599ae0ad9c5f5139baacb976},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{324, 1'b1, 512'h31599cefc10a3c6d549bab5b19bb49d01fad30283d27c8a4905d18cf61e045fffffffff3efa7e2362af0fc827c4bf245dcd58374b350097d26ac996598012290, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00b83f3918b6c5506d648ba3dba36762db593ad4b791456babcc3c1a4966317ae6, 264'h008cd0166047cec89963e9c8ca43b556ac17d0d62177a9bda35e61d0bb16dd471d},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{325, 1'b1, 512'hefe7f8f35a94b65eb3a9299658db8b8256f29f2df969035fe5769c11e85c9b7bffffffff61e57fc3e05c9a1eaf760ce1b13dc6ddc5516048677e1fcd420a6427, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h077858a840230ca21385c4ab4c36cbd3ffaf85656202fba58f1ea995f52ebc4c, 256'h543e5e32a6d2f5c08664ed72175adaa25cdb5d6a754b0cb184e6994ede66c5b9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{326, 1'b1, 512'hc5c3daa9bce3e7422af1de2fdc992b34f5c8ef3fd448b45f2426e1677feaa86aa3ffffffff6e9d87ba471035c9beb5d2c94f3bb0dfb4c48298a8615840c621a6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h538ad8797a397414ac82287c9216e41915c9e3dadbd493a0bbef5cb0dc7935ec, 256'h2c94cfdae7bf76f90b3cc7d19feea4005b387e312ad4116654d63cfbecf2ae1a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{327, 1'b1, 512'he36dcaffe4916e59e41b560c2961fba82290150d1b262323c674311ef6c87564c8aaffffffff573ce47a2b2f25bd4f6468ef2788ede75cd3b7293ad2bdb46617, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ff8bbd1b6441388cb8d562c28ce29fbe51de11502fc825773ded3f0df225b236, 264'h008eccca0148b82fdfb370cdd073aa0634b39cc70d0d5244a7319e4b13791e2c2a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{328, 1'b1, 512'h3f4f00f697d80c258cbcaaeea0f4fa499e0675441a078d32627378ae08c27dc9e8b60bffffffff59976ce86a303743b716e53422d7a17166a185fac1b7722d2f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7c179a010f51d66ec82fe5d5d45bd867b4b236a27be882e627506f7286ed7baa, 256'h5e38c048fb0fbd81c40df3dc16087d9aabeb51a193107499d29d8cf99c388a21},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{329, 1'b1, 512'h21b10973b98ea1dfd2b0d7bfe4adf9d4e8616759177daeef38d7aef0d95d226ec8e1da39ffffffff43f8e40342757a93e72541afd7a58ea2205891c13c72a8e4, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7e0810885b405d54ceb2eb18cae08de2062f61b7ed94ab67eb15e87b64e730ef, 264'h00f511a7919e6e4d70c8d61b831e383f58dea5878a6c8c5f0436ee058dd80a7668},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{330, 1'b1, 512'h3be3c1c0f8b8f6b9c476455ceee9edbf99283f1eab4a28ace9494eae8da166e4aa1d5def8affffffff3d69a06db8c19c0984bdd10df6ede19e4214183d3b0762, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c665d558dd638ef27a28557c3deb8a2f54abf9bd0bfa032c7ec9a514da9a9e9e, 256'h65c9efc355981f91778227eefacf1bb2fedb98657e6cd8674fdd42ae00d619ed},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{331, 1'b1, 512'h14a2049293367e5ace79214bfae58e1007b4977ba9dbd787dd703160651e580fc6de8759ef1affffffff483224ed924c7a2906cccf6b3b39e1af044f2a7047fa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4f06b82aa0d070a004a7fd1135bc3a0bc36fcaeeca35e3edf00f5895394d59ab, 256'h65f71dd7406a17bf19e434a4635479340204dd862a9f2c4653e2fa39b178286c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{332, 1'b1, 512'h745beae01e0b877f882a42a6339b12080d956dfd5fa03fc87f6c99096ae69833fab59c416b092afffffffff5deea8d387d1ecabbcedd6c2334cf7eaa7aa55d84, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h539c8fe5715c3dc893815ec2f00e203b4cd4f8fd36cc5742cc81ced266e02e3b, 264'h00a5964b2d5157624cf42b6726ae23a7d5ef83a5d1f1460bd573d5a15316be5bf2},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{333, 1'b1, 512'hc09dc1025bb9bfa3ef093eb420b7712374f3164db871d4cb44b8ebbeec2d5b415a73427419c5e399ffffffffb45643293f60ae63fb9ff87c56cb45252c8c7c29, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h25f337273591f276849cd855b03d07cbcb205924cda4f62a079591602cc10a8c, 264'h00d7b82c8fb38bbd503d92e5ae9303e8673c6dd0e9389f5af53366bbab851f0470},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{334, 1'b1, 512'h5f9b29b201a8f63acd7387dd71844b5ee67ca50c5a76a2b273a80d167abbdb6727992779f49b848976fffffffff2d0eab3e1c8f8be0d76338c7e8c92174b32c9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00f36018945d24c89678ce2c8cf3cb4f93c38bdad3589891a5baa293744d4daa20, 256'h19ef05878dfc636a4662fd5dd127c908d7948991a324840323c8aef4fc2ff8ac},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{335, 1'b1, 512'ha76f6918ab70eb9171fdaecc8add5917f130dafbb7077543007be1aa2cd3e446114f1fed5989c6275e0fffffffffd7f5a47bd23e9cd47f4572a1d1146b38972f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h43203c89ad43a2bb1910e70ea104347e84764599535d46dabbe547395b1463f4, 264'h00ed3d29c7c506ecc988614b368b38dd5b4f1e330c1b861efca8152a704b9146e5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{336, 1'b1, 512'h1694c34168745c74ab9fe8224e6058e045c73458f7e43e3884e3ed466f716a7406be99e0ef57710a1cac21ffffffffd497d0337e572f1afbc8b6b4f41a873e22, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00c2740bfb3f387df1b564e3ff48835b9e380104716f58c5a43e97bb2c2d84d04a, 264'h00e760ee5d0950b512f6c271cd1a87619b830df83fd40d44b9283539b3aa380019},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{337, 1'b1, 512'h3c28cf3e9527af87b483e6261fe32cee8e67cbc04b983566b27f8419a932186bce21c021eb58c8ecb0b707d9ffffffff035e36909fbfd832447041be74d2ab4d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00ec07ec5378ed131b2dea7ae9776ba536daef2afc38e2556a70b89b9752eb1f71, 264'h00fea25b9e50b1cfa2cf475dbb2245761d5f4585fbbc438d97226c64ff74bff19e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{338, 1'b1, 512'hea6682cf1dadc5f218d6530a15452aaee8857a4318ef3da3cab58358a2e5d0f8fde22dc704453fb8056d224426ffffffff4335e1ab7e6e6c5f3b0a789528694e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e438303ccbbee359c865997e46112b0afd7a647c593429291398f0c432dfb9f0, 264'h008487e07a53da18793f8b527069e620e44587e420245d6ec827bb35cccfae7a47},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{339, 1'b1, 512'h0477828c9cc5710ded82ab21dfa5887f29edfb47548a5a99ff8315da76be5f67922c0a5de1cb7448a3a79b214889ffffffff7dc823ffb5d2fbcda33e63489df0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fc09fa30e89a2ba3d0c4d9d9350e717168c21253371359c0f3cb8c8807bdab56, 256'h5d6c4766bca462cf95b4aeb8f5886b52fc3286642ffee8d0bd7ffd4af7badb4a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{340, 1'b1, 512'h17dfd1c9bfab4afc7d5ac126157041f4c4ca4a04aaf17c45e47857c384fb415e4362041ec3e91609325b7e4c9fb1a3ffffffff9d3efaa9406e392a0dea1ea309, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h4f184fba2be39078385290acb4cc4b3f39b099c3300c762df205c605c6b30e1a, 256'h506481d2018b3a4c0ad558f029c82e0625c833cbbee978bee7b589742ee1e377},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{341, 1'b1, 512'he2fc500440f25769bdfcc82cca36025aa6e5335d8653935dee2cc2a8e8a37c8a886885663c7da8224d2e807f62e1f039ffffffff2aa58c5c932713706022af2a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e9a27533a50eafb09561dc335d67f8e5e53b4fc16b3013f062e581ad027e110e, 256'h7e4150def368f969ace0fc28cac7a3312d6b9af538c412048be1763ea81f3f44},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{342, 1'b1, 512'ha5ce1cdebbed43dea085a592a1ef6c0881660e99434c6f3d6ec24874bb6cc9d56400958f7f95fdc15d3dcc870056263b85ffffffff9f3ace8f83061d0410f802, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00fac24d54387202bff01a91f5504f778c183a0a7930c02af0b618ee64d1b1e438, 264'h00f3a53cb6f96feea45ccadcdf9ac78cd735ec3342163e573d2125caa0d8d507bb},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{343, 1'b1, 512'h6ea638f8043673b9b6a79ff39b5d311774de5f4d697e5251ede52feecabba85d705f25c58b7c2efc844ce598d1428d22e4b3ffffffffc75b0ecb7283d80278f0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h3544590a0f9fa5d43ad4e0a003a8d7db58b8570951657aab3bab732727d1bbc2, 264'h00f257beac10d53e8012ecd236793d280026c5cf1c04aae522019b87e003500ec5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{344, 1'b1, 512'h7cd22c5fec3646707603f858ccd785676b3284b63652913e5581a60e0c262034285489fb945534b7f2578b3e64e7b956bb6586ffffffffc05edada940cffb928, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00bc0726386497c85da8f4055a727b1938e96786b009e6847a080a8aae571b0753, 256'h54b1b15fc7886f09b121af6520d0f4336d259d734713fc3e973cf28368830eff},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{345, 1'b1, 512'hd289f68304c484efc5008425cbf00039a52c7b9d15476d36d58f1515d48a9ec94a850c121249365d7226fb6aad3a82c9eafe994affffffff58e8d36e4237022b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h216f8051f9ceed5b5cc1085f83efd871128cb44b260ac12c486c0ea06c71aa55, 264'h00df90346cb028245a72ac7d8094497f0efb83a7c44ba3b258873127355e3b2edf},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{346, 1'b1, 512'h792eae16afd3069393b20db2ed2e192ffd845b08e10d076d8eafc98744329d6279d31d55ad56a090712fe131358feb130a94bc4a2fffffffff97daeec1130838, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00cb76652e19d6e7a72c9cac35c2ae46178d8c0ff59b06b0cb97c31aad39ec1b09, 256'h5c47b889a29c781540b8783ca24e2acc340178685d7331017e29b4efe92d9fbd},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{347, 1'b1, 512'h51ae80a63d993770d8a5957111af53dabdf3abb9cf9908bc162ded716d3b3c5af2924c076e87c96249a4d7650253ff5112f8a2e7d2aaffffffff66e0e9175efa, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00edfc03190c839528ba2aa0ba3a23b596fcfec1bf2bbf4467f1fd88398cab8ad2, 256'h45b41fa49e0fa7f060ac1ba38ab4d2d5ab5b9fa54ca59285aee09ceedd9865a3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{348, 1'b1, 512'h100c883756f36d7c944d934c08932a99a1c2eb9892cc39a13a80b22aadc526ad755265f9ebbc8d0c1ccd31240299c71604332ff56592b7fffffffff1224308a3, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00e7631f03d9dfddc64cfd2a971523def68cb9f8a64e07eb2235c7250adc36480b, 264'h00a004cbac3e04056c7e65fdb48be051e9a52ab427c826c84e2cb2229252983663},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{349, 1'b1, 512'hf4272253af2b51df321249280f3f3e62fb1e4a4a556f88bf3d5ae20ac5cc3e035e7b2141f9139b2f21d431068b8d5d96fcaad0f106289298ffffffff51777f01, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h15e36a42515118021f6f5372ecbff90755d8ae77f9dd683972d2f26aa6716451, 264'h008d1cd988ba0a1bd919d2f9b5c8a3517eb59ef776caecdf2b5ac2f7a721858315},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{350, 1'b1, 512'h8bfa5531067a5cbc9bf002be2397bd10dd183d7ae47a02c0d0a7d87e1f94af93ea7365b711cfa611750ac963de0551c900dbad9cd8071b503afffffffffe6b6f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6daacbc1125cb3690e43e16b414077c0dd274b96ed61892bad5a519274f01b23, 264'h00d044965811b4050c7a85021e8827635cf9f46260fc33bb7cb56b1b37180c4220},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{351, 1'b1, 512'h8a5409853b325b917b8a2aa1eb394767bb07fa82af11357e777f7404e0955bc9bb9cc5a918475c52df4772a1207e3ee4f3e3d3c8e68e84e10477ffffffffd35f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h37e50775ee06024d596ed49824b1e6a49efae25c7dce8181de33f93ce34ac3ce, 256'h616a3e9d1fed086138f6feef6532647c02bd324ba4a8bfea20640d22f5494429},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{352, 1'b1, 512'h8e38a571ec826b9af00de0c523b6e073aaf9380cc64fbc86755f33f065361d8963ea2c42796ac7516f53d689e1da364bb7caf6b22a5fee81410646ffffffff7f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00d5b64cdf82e354ba6a01772f7d38e8d46a729b808aaed73616ed41a9afc83db7, 264'h00b5c456c91254e57013228c9724bb7f97aaf18e1bfd4c99d3ca9eaa8214382a10},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{353, 1'b1, 512'h0f3ad12803aaf9bc615745a47da85dd90bff191d3e9441cc2cc96bf8c01f5e514b256685e3e48f01a98a5f27d20cd1c317a6f816ca8611fbc8891236ffffffff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 264'h00915779b90ae6f6c1fb82c198c9f0719ce2ea37be0f261e36585ec89adaedd2b6, 256'h7d05e7794ac57578790808c0ac52ca3a51d1399f1a4c7173a7ed19867732b3d9},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{354, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h097a04ee03a13c511d939e8bbe1471c57a71020e168e2689c69a5625686e24ad, 256'h40d24d52f3701ac8da959560c36ed0750a1cf031b728a9134e2b71ed3ddef889},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{355, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h12c90a5debd88d42686b84227dbc755351b78e7c6cb86c0b22536f394603646e, 264'h00d03d965851bc41bb089499c51987b899a8353d997e040fdd35290a2627f0a3ab, 136'h014551231950b75fc4402da1722fc9baeb, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=136b(17B), s=264b(33B)
  '{356, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h12c90a5debd88d42686b84227dbc755351b78e7c6cb86c0b22536f394603646e, 264'h00d03d965851bc41bb089499c51987b899a8353d997e040fdd35290a2627f0a3ab, 264'h00fffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2c, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{357, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00913ed043022ee590f59e44f519e5cfd9d6f1b84a50fb417e9ad06683c6afa194, 264'h00b68fb80d6ef261b5a63b57f871d2ea7224319f5fa3ed3dd77f1012dba19d0395, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413f, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{358, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h644cc54e84467213fafe2a4451dba550f3ea76ea9970bd6251fc7783a420d8b5, 256'h1cd9439155ec45d5634677c281154bbdf99fe44051dcec322053ca69ea88297c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3e9a7582886089c62fb840cf3b83061cd1cff3ae4341808bb5bdee6191174177},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{359, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h0a11d42154bd2de10ca92321fb6b3e638ee8b5a7fb4fb5f501b44515cf60e8c9, 256'h06ccaab8748cd38ece73ddc975bc307e7de172357e14cd96a94bb3461d32d50e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h24238e70b431b1a64efdf9032669939d4b77f249503fc6905feb7540dea3e6d2},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{360, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h009fa2c32bb349846acb5af14e1c67acfdd8963ed251c4b5783cad4bcdd0fd505d, 256'h6f724937217d1e5483920405cf1b20200797521c464a2355fdde5306f2a9e448, 8'h01, 8'h01},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{361, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h60eace95001201cf4c83b580fb698bb6abf446e5c56ff945eb5769b1a477b550, 256'h69f5354a77fe2d601528f126c9a6858deeddb9e5ec408356d05ed5c80d62b8e1, 8'h01, 8'h02},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{362, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00f1a57d9346842310975ed356672a48a06a70b5efbc0c23287c9b9952ec955b33, 256'h0091aee1224ecd69791856c521b12df172b45a5ce247e6dcaca7349684278f23, 8'h01, 8'h03},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{363, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00f1a57d9346842310975ed356672a48a06a70b5efbc0c23287c9b9952ec955b33, 256'h0091aee1224ecd69791856c521b12df172b45a5ce247e6dcaca7349684278f23, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 8'h03},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=8b(1B)
  '{364, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00968a493f279c0f8ea9f2446e361ee5b9757039d57a8003e6fd731d4dc6a2d2ca, 256'h6784c5484fe797c830aa49a72cf85375523228393b730b20b04a192032af4d29, 8'h01, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd04917c8},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=8b(1B), s=264b(33B)
  '{365, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b3c7fbdf1d7472f7bd578757762c8ebc922ff063b0ae9c3aa9cd81600abea76c, 256'h038eeb3852b836c0649fd82fe5d1d02c3d0dbb30fbcd7fe41866ebc3bd927c69, 16'h0101, 264'h00c58b162c58b162c58b162c58b162c58a1b242973853e16db75c8a1a71da4d39d},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=16b(2B), s=264b(33B)
  '{366, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h759fdd1a64c000188b87eb0ddd291a50358fca2b0a5b92f027573845dc40b27a, 256'h12ec1b2892ef46700f13cff8eb88f40076cc811478b008f5aabee4a74b4546f1, 56'h2d9b4d347952cc, 264'h00fcbc5103d0da267477d1791461cf2aa44bf9d43198f79507bd8779d69a13108e},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=56b(7B), s=264b(33B)
  '{367, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4882825a892d30267264e300e868ab5d4b0ffc9ef3c2cb6e90d61d238daed856, 264'h00e4c8248a189eb36d83740f5928cb802fb9c50b5a18c9196344a0c2cb74416423, 104'h1033e67e37b32b445580bf4efc, 264'h00906f906f906f906f906f906f906f906ed8e426f7b1968c35a204236a579723d2},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=104b(13B), s=264b(33B)
  '{368, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00c4d1b1fdf274cf83f3395a70a36c94f7c51f1a31e99514b4ef10ba1304756caf, 256'h4eaf435b20dd76d6ef447869503da9b28f0ea08edf287424d44aa04b254c1736, 16'h0101, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=16b(2B), s=256b(32B)
  '{369, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h3376df7376d5e651d45b8ec2e5ff9d891c6fdd6dbbb52b046e6b5ac4c9facedf, 256'h76cf27f9fcb65403b1f585a2dafe26b43ebd622baccde699d81c9be98df9f4df, 104'h062522bbd3ecbe7c39e93e7c26, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=104b(13B), s=256b(32B)
  '{370, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h5077fdd202fdb4194b05491b6c053fff8760697531fc5227879e9cbec3309585, 264'h00d0b5cffb3e0fdfb1c06e6d11a1182752730cfe439f7a4f8a49b9c2924f49ec14, 264'h00fffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd03640c1, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{371, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1b1f773b472dac5e1adf94e69d865b404d2cc92cff7bb66cf2197978f6c45d08, 264'h00a9725791c5f33787977a9ddfa69296be998a968c51ec7f1c5447793bc56286b3, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h01},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{372, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1b1f773b472dac5e1adf94e69d865b404d2cc92cff7bb66cf2197978f6c45d08, 264'h00a9725791c5f33787977a9ddfa69296be998a968c51ec7f1c5447793bc56286b3, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 8'h00},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=8b(1B)
  '{373, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h2f20bc2232b4ba9d75fea6a92bc827d91c5a8f5c887f4e304d76656ba15999ea, 256'h5f83242efbd57dd16dbd3de0915bdb2ddec201d2f749b13fc22c223a2644dcdc, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{374, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h009e009cd0a1a7d0c51765169c468e62e56fc4f3ff02e8666c55483419a2560032, 264'h00cd36d713acd504598ff3b4f58046a4690f550bd60ef4c823c5c581c6b899315e, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{375, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00af58a6ecc8254b9b831ae0441c13990802c3d68c301d43634c71f1974c09e704, 264'h00d920612d82f32fca436c5c5097505271494875402731d03dba942b355306c783, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a1},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{376, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4a7217cabc95b496f3f4e12d54e9def7651b866be69d3695cd77ad2e3a3f13d1, 264'h00d0fa71bf21d2c00b1ff4cc76b53a9c5c2a8a8b6b4c2ec88b99ee537ac6262b3d, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{377, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h00a42e277ce657fb3dd07e135a3cb9b0a75a30bd8b64911606ee68371e561244, 256'h67cf22e26a7009045b73ff19cd79851cceaad9ae72ef2d043d75365245befa06, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 264'h00bc07ff041506dc73a75086a43252fb4270e157da75fb6cb92a9f07dcad153ec0},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{378, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h008520b9502f9a5ed753f09a5282cad721f5ebfb3db4142d667c6279869e76bcf1, 256'h678e9bbd04a51460afc40a3e0cb7b0f8b8add89b2979758a5a1ffeb4584ee49e, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{379, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b5deca0fe0296905aac27e3604a95a0a2ecbee9fc453d2e1164632964454d0c9, 256'h4f9e4e85a143ee677d40919c71014e8cabf4d9db7442fe4b96298f99f90ca67f, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 264'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa9d1c9e899ca306ad27fe1945de0242b89},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{380, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h5dcb2767dc851e20911ed7be39dd87ba81c7a6d10255dfb825f241486f98ae10, 264'h00f8a9ef736b3e11d7d54a0e086902fb477246ec8c57de65d336570b65f65e0d83, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6bfd55a94e530bd972e52873ef39ac3e56d420a64d874694c701e714511d1696},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{381, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00c8e144c853a7e1a6f5bbabe7ef91ef5b152113210d44fd58d3cb6185184e168a, 264'h00ac40fb3618882193fc6d113760e476465df49067480a0a7cffe686515b3391a8, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00b494bd67c209a5adb1c9a09337e2629b03f8a924be53c542478e5864ed2622ad},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{382, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h7ffe185a23eb5b736704387e6357628a65984985773b4473cf9ef560b3fa5051, 256'h4740cb1217f1ad2b5910d7f74906602b1f9550b3d11cff705b358c3bcbf72c3d, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00aad4e2b69a9f378dae7873b40f7c15cb4565fcc8cbc0ec55b0bd3fe9d8626b2c},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{383, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h008a858226155e34dbb7e5dac7f13127c81c6ce8c9d891918c67c8738d7e4b46e9, 256'h6c1386e84c612312de53e9e4af34d9bd57f93d9a06b855b6e0b06ad4137ff57c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h73fec4995e9d3140bc07ff041506dc7313e95389fb599d22f24039392a4014d3},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{384, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00aec0be729b02f266c542d139a3e04110c933e8eca1008e8dba38d75e7f8fab53, 256'h2cd688d924b456848bd5c651444c67a9399fdfb5b5b9693162c1728bfadc1046, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00ec4995e9d3140bc07ff041506dc73a73dc25f4257a911e310e38744b482a5a01},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{385, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h01ed4b5f941f443b31a7e2583ea165551d1815b54740deb12e9fdeff32e23061, 264'h0084385ca448cc5dd71139bda3ab42d0b6e44d719e52fff64d971876efa9109fb2, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00d8932bd3a6281780ffe082a0db8e74e8fd9d0b6445d99c265c9e8a09c01e72c1},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{386, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h59c427cb6525eab511a06e03e00cf2aab4abc587c2601534338a50bc25701a70, 256'h3e4eb388b453cbaea594d6b5c14a519ac3fda770c53580beefc68f09200d55ff, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5e9d3140bc07ff041506dc73a75086a3ba176f06c2b6e37363e2ce1c141f3c27},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{387, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h04acbbcd23cf2ec819fd297ab2cb5407ede6319518651a391e941cc800356833, 256'h1206dd00df23bc8ce0b85a018c4b34e9c3b41b4ef59c71492fa62d134772f97e, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00fd6dc71a71f1d50d1bbd976af4357be4dd2fe850707c431fd376e53d176c6b62},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{388, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00ccacbc626fd6ea31175815cff958ca1637323877d3bdf09896b527bf4e255e85, 256'h71f8a27e6309bd9b9b15d78d5270012ad2ed15a7fffe024fc0eca63fb6ac2f8d, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h7ee75ad2a5801c54722eb7d95ba67febcfc399b956b7b682fe89638de3690bf1},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{389, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00ccc30b65cad3dd1d793b6db80f57b2e1237973e4264c3d9bbc2551ec68a0b7be, 256'h75ff6d1f4f535a131aa573f6e2d6912c397154933750417d28e46524392592de, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00f533776f11c47ed0a7b5e25ace7a3b921866733c7454b2c678b8943dfb4cf232},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{390, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00cc9349aca0cbd0b2df0deecd88ed39e6d8c7c3d7b422fd5d92431baf7225fcc0, 264'h00ed494be698d6f3850be277c268792400f396025cfa95cf56018bcbc243e512eb, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00e8dbffee01807d75f9aa52c295e15b15f138439e7a195a40709b1abf511dbc6a},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{391, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 248'h0e7c30d2f259f7c13f194320e43905d0ead7277e283e8918437c10f9d052b0, 256'h2b39b66dbba2b1cf5dac1b41d2dec6f1fb08bdd14d420d703986f63aedeb5c47, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00ca01552b58d67a13468d6bc6086329df8f44cc938884fcf15c516b02a7a7b5f6},  // lens: hash=512b(64B), x=248b(31B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{392, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h008fa298c00ac93f7c36892c5299005a0f6843f9cf0669fdbb7d6d81e0341803ed, 256'h4cab33cc2821b2da849f90ef20dc1eb896fc67161440b3c52c0b1e88627e508c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h009402aa56b1acf4268d1ad78c10c653c063dabc4061c159a6f8d077787f192aab},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{393, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h6fbf608a83e37ec26b37da033e069816680b770ba766fb8c44fce003960562f1, 256'h045f268ccc5e0949213f7f2f1fa57cfead04625ec3ccfc9c333596e487b2056f, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5e03ff820a836e39d3a8435219297da13870abed3afdb65c954f83ee568a9f60},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{394, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00c4dd547ad750174179bac8b8ce27481c58b81347776220a1b52ada13d65c8124, 264'h00f9c2ef3b5b4957cf69d3a139891682363c040610f200f4c318e59aa68f298af0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h556a715b4d4f9bc6d73c39da07be0ae5a2b2fe6465e0762ad85e9ff4ec313596},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{395, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 248'h055d79fb26286bb6289a7983a2b23bf5c30cc3d70363b559adf5548af991f8, 264'h00cae8b1b0ace32fd74a86ee1a671cc36c052a4796eae323be32e02ce9a0fb6227, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00d55555555555555555555555555555547c74934474db157d2a8c3f088aced62a},  // lens: hash=512b(64B), x=248b(31B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{396, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h0db51c74d34e41baba67c13a60af404ee82d8f1b0386b09696ee1e6ea1327b86, 256'h413886c4623fc222a6950c3c3a09f3fd867a566bfd345e06b09ec6c5c2e4a192, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00c1777c8853938e536213c02464a936000ba1e21c0fc62075d46c624e23b52f31},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{397, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00bc2f7bc74cb3bc7e797b06cc3e649bf3407d1a55b4eaaddd28d3dcfaff2c3737, 264'h00a23bb364e16ac79398c013ce29a22e762c0d6067aaefda958474aad194a92e8a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h30bbb794db588363b40679f6c182a50d3ce9679acdd3ffbe36d7813dacbdc818},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{398, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00d7edc7c645efff6af8821aea5b7f969f56ef6e615862b08fba3eaf0111c06f67, 264'h00e47fd0da61682adcc405f329148bf1c35b89cb5ec5a9ed0d98a410e261a6b41a, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2c37fd995622c4fb7fffffffffffffffc7cee745110cb45ab558ed7c90c15a2f},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{399, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h6bfd7ad01b5dcfb04de464083d3ca7ef5054506111df92ef02ff7690d9a6ec93, 256'h06c469fe4c5a1e04f114e193b4bb197de2c8e35089037e5a20275bcf67d9bf73, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h7fd995622c4fb7ffffffffffffffffff5d883ffab5b32652ccdcaa290fccb97d},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{400, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h008a9076c923021d5c5ef85894176ebb5c3a74aba75b3944c96f17debc2173ba99, 264'h00e5601d115bf08d37ae115c4d186bc21127bbfb21d0629bde27a16e9ed721b740, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00ffb32ac4589f6ffffffffffffffffffebb107ff56b664ca599b954521f9972fa},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{401, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h0fec6a85e077ef4240b98c62ab3b93e2cebcad0ae9617f7b0471504db1f45a65, 256'h245a5fd0ad7a6d854125ed76d4787f77cc1983eca8c6ba8c019523a088c4d0f3, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5622c4fb7fffffffffffffffffffffff928a8f1c7ac7bec1808b9f61c01ec327},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{402, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00d3ab94d8704fb51774dcc3838ad9703071e0851de9b2d6ca74ccd79b85558191, 256'h4e4979b67f377419e5a9d4f03012b7e75656556f23756d4dbee145834c8279ef, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h44104104104104104104104104104103b87853fd3b7d3f8e175125b4382f25ed},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{403, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h49e13cd44c8b8350a5eaca2181bf96db120b768bde8800f379f43e9198333c75, 256'h030ad9fb4b0b233bdc10ca0dc4c2134b18b691e46c7151e3573aa2b62891e69d, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2739ce739ce739ce739ce739ce739ce705560298d1f2f08dc419ac273a5b54d9},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{404, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4574fd94ad03828588cb0bc2d434842ee093efe639015cc107d1ea3710f2112d, 256'h1786d6ef1d411cbd1af5b5ee8845993e738fb64519b4329d04be21f7902a1c1d, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00b777777777777777777777777777777688e6a1fe808a97a348671222ff16b863},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{405, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00ee824d818768f13fa0eb908e396ea1c56b11774ce69d01e563aa36bb41d6371c, 264'h00990291ce2abc55bb6682d502ae0129e7c57e146e96d44757daaa1f94c93e0b17, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6492492492492492492492492492492406dd3a19b8d5fb875235963c593bd2d3},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{406, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h4825ee46b2d21564726a32a922f5e3f2da6098f780e1f15c6bf1640669c41fe7, 256'h292c066a24f0f450c2603f1837210898f8e80fa384aaf077eb5c7e87c6b26976, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00955555555555555555555555555555547c74934474db157d2a8c3f088aced62c},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{407, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h41348e7ac18eb1f4852801467bb0a0e36209321a8af4b410fd06f070a81f5de6, 256'h03b5594f1a5a79d23089e49e3e379f2a6cb14f92301c6999e510b8c8dc37fb4b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa3e3a49a23a6d8abe95461f8445676b17},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{408, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h753c74e5a36e1a4b61be7787202c98e05841fea2b0392b6ab69ee2e8a747e2b6, 256'h18971da1c85825c1d8141886115d27cb2add86545e6971bb835a2f452cde1e52, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 264'h00bffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364143},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=264b(33B)
  '{409, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h49c0254724576b0949827ce46240d90cb4075cd1978a416495a455f06a895504, 264'h00df7d64c35853353bd4d905da6adb88f26e62a5f20b3cd6382adf2c5a42d85053, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h185ddbca6dac41b1da033cfb60c152869e74b3cd66e9ffdf1b6bc09ed65ee40c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{410, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b05e98e84e2c19743c1dcf4e0ddf0bb1f32854033de63fcf3e605fbb2ed94cb1, 264'h00871d7415d5f6c57c840678f7e1a1c1e323519a4647fb3f6f52abb4647b9b6d70, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 256'h6fd848306e968e3ac1f6e443577c47a3c20bf0d01a5dc39c78c2c69d681850f4},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{411, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00b05e98e84e2c19743c1dcf4e0ddf0bb1f32854033de63fcf3e605fbb2ed94cb1, 256'h78e28bea2a093a837bf987081e5e3e1cdcae65b9b804c090ad544b9a84648ebf, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 256'h6fd848306e968e3ac1f6e443577c47a3c20bf0d01a5dc39c78c2c69d681850f4},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{412, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00a49f9ebc082c064d61c0eab5f8bf23207b06e3a689dfc4fa2896ed114d1a88ab, 256'h55783a6baf9401977d117ccb748c0d5c24a5d3bd2133d62c74de2be7cc7d9d40, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0, 256'h33333333333333333333333333333332f222f8faefdb533f265d461c29a47373},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{413, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00f9567a431b716388428510393b37feefd3afcfc6dc3881f623c0a0995e461ec3, 264'h00fba2f910ced19f8e789b158390a295e636c588c622d54f8feffbd2852e2911a9, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{414, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h26095ef93b10bf50fe283f4c99136fb81fa297814f09977e8e38a3bfb837f61b, 264'h00af8d7cfc46c1928624f201ed14a70701bc5531bff4e2e578d5c92dabddbc7580, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 264'h00b6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{415, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h7a4b58ee76d461a1c3cde68400a0bbeeab346ee69315bed63f1700c66cf5e6cc, 264'h00a642ae4078bb6bbbb76028977882e9c8374f267a2ced131029ae89560ce29825, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 264'h0099999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{416, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00f2a111eb24c9d280d9a66e4ff18681d222dd6a1828ebc4528f2bebe3e25228a1, 264'h00a0699bcec507fd0ec83da541a5a6143e2e68e4af72fcdcc8a2aea2b17478cc8a, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{417, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00e50054b3e4a4d1fef988e5a5e830155abc293fea3598af4c5ddaa10acd111274, 264'h00eb710d1834568cb379a1d1f3d691a8c0dc19f901fe3225c2b6691df5ef5333fe, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{418, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00edc17cd4ca6f9988fda5af4042e3f9eb42d0f7b6a1c0156e1a2af566b7810354, 264'h008a5d357777b306e96405f12e2617c1b29e8d574e5f6d66d1bc8ff7ea7c4b683c, 264'h00c6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{419, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h6d267c10d2315b42dbaf34c97c3c0d331fabacaf6021df4dc85b3e9e63dc0798, 264'h00ed154b11fa3a5ed952c14d8a2dd242de2b6cce3c22df42cd97de30054a19555e, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{420, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00c24bf7a984c96ece10077a9def38cbd0d898abd555f1668e06c27cabc00f6f67, 264'h009f69b238e1f95e99e5b558e0036273ebd6c36d12b4515348b85a21f6283f5016, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=512b(64B), x=264b(33B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{421, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h1cd26d668807c815ed3f532c1db81ac473fb368f0f7ef1aff2592ea6fa6c4624, 264'h00a229b9ab5746cfbc47280c019a4248545354ca20880ff41cac2e252bc9b49704, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h0099999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{422, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 264'h00fc780777a3289af663fa02b1c262a8373b84614e659c1ab46942f1e058926ff8, 256'h2196c6bcae0b2798298d463be5c87924343d7f103a27131e0c7f4d60d2b5da8c, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{423, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h5e25e2ee8af5ef8a3e0908341f9884501fb58a2fd234b1db6f22d561025524f4, 256'h491d97a7793c9d9a1f35bb35f12121b9dbe075d8501cbd4db6697e3e0ad98bc0, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{424, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h3ddf2920607df596da90123ea5674958054c8ed7758661b813f1aa30f19778b0, 256'h707243e1a7bcc264b54289832e950c27563856241b79c243d0fc54f7ad24bc25, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{425, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 256'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{426, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 264'h00bc07ff041506dc73a75086a43252fb4270e157da75fb6cb92a9f07dcad153ec0, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=256b(32B), r=264b(33B), s=256b(32B)
  '{427, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 256'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{428, 1'b0, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 264'h00bc07ff041506dc73a75086a43252fb4270e157da75fb6cb92a9f07dcad153ec0, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{429, 1'b1, 512'hcf83e1357eefb8bdf1542850d66d8007d620e4050b5715dc83f4a921d36ce9ce47d0d13c5d85f2b0ff8318d2877eec2f63b931bd47417a81a538327af927da3e, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h6632473c909425b6fa37095398e2538daab8552440320f9fe190dba8f672796b, 264'h00a8c3aacce9ffe4bc17c0530738f1386f9d9579f029ff3a7791b16e98422265e3},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{430, 1'b1, 512'hdc5e71048a56da7aa1bf5fad1ae227446663488d8a531d490c4b5efa048ca4651acd9a196d9b13ee2a1c74ad440bdd88f6a34a02fbfadac2f7ce869e64486558, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h465b0fb05c14cd4ddef23e13acbe5f2337c45ea3816536670cfa7f2ab9090619, 248'h5e525e837c406cf8944383e20bcee32112d8da5b42b40f88415098f722aa89},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=248b(31B)
  '{431, 1'b1, 512'h43f800fbeaf9238c58af795bcdad04bc49cd850c394d3382953356b023210281757b30e19218a37cbd612086fbc158caa8b4e1acb2ec00837e5d941f342fb3cc, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h7b1553e4d650c71fd49aa36ceed56f0438b0065e1b234445134bf7c83231ca9d, 264'h00e369a20fa6434bd138b092885a89e53a3f0b6bdcc5d2653e136c54070081dc5a},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{432, 1'b1, 512'hd296b892b3a7964bd0cc882fc7c0be948b6bbd8eb1eff8c13942fcaabf1f38772dd56ba4d8ecd0b626ff5cef1cd045a1b0a76910396f3c7430b215a85950e9c3, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 264'h00c7ba1c73bdc4364f6c7c61ab1fecc0547f8d6fcbeb251f734964407536353f32, 256'h7b3a6fb2fe60f8861e9e0955663f5703a17f5ecc3a5b5140eb87eaf35a3a5090},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{433, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h2b9c9f85596fed708b3af80393b27edfd0b5ae2f0074270a56362f5f9f62b4e1, 256'h2fae837503ba2c1d4c945e0913949ef094ce0b8086359bbb5dba4a12707c5600},  // lens: hash=512b(64B), x=256b(32B), y=232b(29B), r=256b(32B), s=256b(32B)
  '{434, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h5cd765209021d8c1a8aef4ff61d6fa6e7993bf9fea0b93609eea130de536fccc, 256'h4f10c7989587fe3019e36d85aa024bf20db6737c4f28900c1c9662f2782143e0},  // lens: hash=512b(64B), x=256b(32B), y=232b(29B), r=256b(32B), s=256b(32B)
  '{435, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h4c1a59b1e578d76f1595e13b557057559f26ab559ec1df3f45ec98b90fa526ce, 264'h00c6872f094bdb3f82e31f93ad65357e2daafe66f304af197089ef0dc94ff90624},  // lens: hash=512b(64B), x=256b(32B), y=232b(29B), r=256b(32B), s=264b(33B)
  '{436, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 264'h00a35d1400d4cc7a8f617b721faee7118a74103c4630dec5aa47e097951dafc1a7, 264'h00958221023024e97ef6df35a22e820c7bc5e16299f3f12e9d9b1b727c46d795e6},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{437, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h7fb733ed73c72fc4f4cf065e370c730301316ff4e9c6a8a701170f604c2d70b7, 256'h7ca9ca985d3df48978b3a2f9c0bb8a58b216c795e687f74623a3321448bfa73c},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{438, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 264'h0095ae4df2fba8524e1151cb9a9c5c1ec1357a663722a18329303d86a58e704754, 256'h591ea644b1dc6f4c7cd5d7d939397f84d9e077100760f0816ae5b22ae6a74203},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{439, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h717925f0dd5cf45e746e87f79c9ea97d11eb01444052c270aeccef56c2e95828, 256'h785787b664137080383d2fc500459fa713258205fdae97b3240fb64bb638a657},  // lens: hash=512b(64B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{440, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 264'h008adfdeae3b586315d06183610d271fc423cc789908b8f5dc563253a3c782510a, 264'h008137bedbb4e60da26041b351f72a6bc3b7741f745743f0733b40b7fc56febd04},  // lens: hash=512b(64B), x=232b(29B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{441, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 264'h0092ded14e19b94d17c79b063a034b122ce3b93a2502f2f223fad3461abf631632, 256'h52ff8ad14ba3657242e29440d01cab36ebb6033ee36021dc8d9b38f0808a90bc},  // lens: hash=512b(64B), x=232b(29B), y=264b(33B), r=264b(33B), s=256b(32B)
  '{442, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 264'h00d48373483e0fa2f11cfdfaea6f1de59e6861e9e87c4f6446602ba0125ab7de46, 264'h009d753bba3a7be08aab456e93a6500d4781795ed59af8bd6d6133129abef1ad98},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{443, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 264'h00f11473117b66e5d84a2ecd0f8b7ec4a2cc2aee89ae022020235777305142f498, 264'h00fe5ce43ced28f3f69f65e810678afefd2bdeefb051280ad2880157fda28b2ab1},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
  '{444, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'h3c9f5bdde7310b5696c93c86203fc97e11a70739e20c71c9e722308d45a59e6c, 264'h00c09efb9a045a47cce799b768890bb17833a0210d869a36be1da33f2585477c32},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=264b(33B)
  '{445, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'h6953442c487f240487d2af81f9825c894b1fc2534321fa012db8248be20a4b06, 256'h56927395d64ce4d690caa98944c2ddebc312f57f439d37236ea63cc1de098718},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{446, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 264'h00fb39aa5f36ceca6e68d1932e811598c412892734dade389fd9e8ba94c5c7a251, 264'h00fdddf0c3db66c7c46608ac98431f0ee8ebb1e27ba501937789ebcd0f7ac26ecc},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=264b(33B), s=264b(33B)
  '{447, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'h44fef6017638fd5bda17dfce346b0311b5e369bfb68aa85d5e970786b8e6644b, 256'h720b3a52fe44be6028759f0f1a6fd7020ff6792cd4ece98dffd0d97d3b726091},  // lens: hash=512b(64B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{448, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h304babc41346e6205cf03e2d0b26e4b222dce8227402d001ba233efa69c91234, 248'h65add3279f51b2417fb0a13b0f06404199caac3430385513ee49f67d8e8cdf},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=248b(31B)
  '{449, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h23868700b71fbafcaa73960faf922ee0458ef69e01fb060b2f9a80d992fe114c, 256'h6ec1526bd56f6eebf10463bd9210d62510b95166365e10a7b7abfc4d584ca338},  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{450, 1'b1, 512'h4fb472dfc43def7a46ad442c58ac532f89e0c8a96f23b672f5fd637652eab158d4d589444ef7530a34e6626b40830b4e1ec5364611ae31c599bffa958e8b4c4e, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 264'h00dd60d7cf83a08208637212b65d079fb658d8ef1b8438d9c58f4122b0cd14ac49, 264'h00f1d762516f4d6c3e6a98dd31dc3869dc7cf35944f33b35c6a17fe632d2b18cd5}  // lens: hash=512b(64B), x=256b(32B), y=264b(33B), r=264b(33B), s=264b(33B)
};
`endif // WYCHERPROOF_SECP256K1_SHA512_SV
