`ifndef WYCHERPROOF_SECP160R2_SHA256_SV
`define WYCHERPROOF_SECP160R2_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp160r2_sha256;

localparam int TEST_VECTORS_SECP160R2_SHA256_NUM = 230;

ecdsa_vector_secp160r2_sha256 test_vectors_secp160r2_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'h00c85b8de817a9a998acf135a918c146c7ebde2b3e},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{95, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 176'h0af8cf160e6cdee66be28cc2e341d85210f931d00000, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=176b(22B), s=160b(20B)
  '{96, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 176'h37a47217e8565667530eff75cec5615107c3762d0000},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=176b(22B)
  '{100, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 176'h0af8cf160e6cdee66be28cc2e341d85210f931d00500, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=176b(22B), s=160b(20B)
  '{101, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 176'h37a47217e8565667530eff75cec5615107c3762d0500},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=176b(22B)
  '{116, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=0b(0B), s=160b(20B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=0b(0B)
  '{120, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h08f8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h35a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f93150, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c376ad},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 152'h0af8cf160e6cdee66be28cc2e341d85210f931, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=152b(19B), s=160b(20B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 152'hf8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=152b(19B), s=160b(20B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 152'h37a47217e8565667530eff75cec5615107c376},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=152b(19B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 152'ha47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=152b(19B)
  '{128, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 32936'h0af8cf160e6cdee66be28cc2e341d85210f931d00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=32936b(4117B), s=160b(20B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 32936'h37a47217e8565667530eff75cec5615107c3762d0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=32936b(4117B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'hff0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{131, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'hff37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=8b(1B)
  '{136, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h010af8cf160e6cdee66be2c1e1cac8806b049ad33b, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'hff0af8cf160e6cdee66be257a3fbbb30391d579065, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{138, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'hf50730e9f1932119941d733d1cbe27adef06ce30, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00f50730e9f1932119941da85c0444cfc6e2a86f9b, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{140, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'hfef50730e9f1932119941d3e1e35377f94fb652cc5, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{141, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h020af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{142, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'hfe0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{143, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h01f50730e9f1932119941d733d1cbe27adef06ce30, 160'h37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'h0137a47217e8565667530f3494b64c0969fb651798},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'hff37a47217e8565667530eca56e73eb9381421d4c2},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 160'hc85b8de817a9a998acf1008a313a9eaef83c89d3},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'hfec85b8de817a9a998acf0cb6b49b3f696049ae868},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'h0237a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'hfe37a47217e8565667530eff75cec5615107c3762d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0af8cf160e6cdee66be28cc2e341d85210f931d0, 168'h01c85b8de817a9a998acf1008a313a9eaef83c89d3},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{153, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{157, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{158, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h00, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{163, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{167, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{168, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'h01, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{176, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{177, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{178, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 8'hff, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{182, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{183, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{184, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{187, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{188, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16b, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{192, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{193, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{194, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{195, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{196, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{197, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{198, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16a, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{201, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{202, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{203, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{204, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{205, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{206, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{207, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{208, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0100000000000000000000351ee786a818f3a1a16c, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{211, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{212, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{213, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{214, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{215, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{216, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{217, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{218, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{221, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{222, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{223, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{224, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h0100000000000000000000351ee786a818f3a1a16b},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{225, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h0100000000000000000000351ee786a818f3a1a16a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{226, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h0100000000000000000000351ee786a818f3a1a16c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{227, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{228, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{240, 1'b1, 256'h85ea0bd8290e936b523066a9a85c32fd33a50dea0855f5d0c4e029a4a9ae7365, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h7798282cd94abd9bb74be4191d4c48755b515f27, 168'h009363c32313f924ac79172f58465baebe8136ce22},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{241, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0084796df79b732a372f94e18e50a58e5f8ded936e, 168'h008fc1eccd24f4385a611d6aa7ae3bf185e541c547},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{242, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00fbd482bd1f9c1fb279cc08f2ef8fdda23616ddd5, 160'h3a0f477b82bb13ad5c3d44bdf2835f2c434897e4},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{243, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h39b0c99df627abb063501b93bc0ec2f9fe1abac9, 160'h01e957fe1c54b5ba221f79b64fc2763fffa80524},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{244, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h2ab314be8a53a6af98e60e9378ad5194a6306629, 160'h60101c49dbbcf678851f678562bb99b0e983d011},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{245, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00a67d8de97700cff561f4f089ee06a07f11ae497f, 160'h675a4ee3a50a32f1d7fd5503b820ddeb3b1c84aa},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{246, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00aec171c491b59627dc9c50b5c7bfaed71b5d8cb4, 168'h00d388a785cffb83e294cf74210b31eaa48e9e7081},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{247, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h1ecc9059b760b9561bfd933956241a0e33551f9c, 168'h00c0ee636c93c6f3c48f2705226aa633ff58831796},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{248, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h53f4103b4ff5f2b04e60409b712b24e52d446bee, 160'h5a0a9c4e5ed87323e7a2f8964cdd05aaca8623f5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{249, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h623a961ae133e8fcc433d41afbc7d479bbacf5a7, 160'h120f4662c44fd860a09057d016ea22f59c9ea48a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{250, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00f73cc481f89915c1c5afa325f669d13c99776a8d, 168'h008a3a09961127584ced19d4c1e1783b60a8199a0f},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{251, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00b3f652bc6bd17fbf0776179c1ae506a2bbe177ce, 168'h00ca8abc2878a8cd46bcbc5a4dba835d27821eae26},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{252, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h2381092416200a5a4d79761a6e5968ce29507e88, 168'h00abb04b04d8e5d606e5b0aef01833df967e04bee5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{253, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0b1f411f5693fb1dfec23bc48e415c83101c9275, 168'h00ed771f55741c53446b3ddcbdcce143774a1de7d5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{254, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00846052d0a5a8e970c22600710a030739d6636545, 168'h009d8ac70e6a74cf2433291a96134339fba6c08d38},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{255, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h55a270df082a4d6183a4b6ff10a737e02c48b4b8, 160'h5026129206b77d6b0de92147deb0d0ae7c2260fd},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{256, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h6d84f406773166c41bb442f5af04ab9858df5604, 160'h6aa89196cf9bfe8dbcda618438dc717c8fdc0bc0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{257, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h015667f4c09576876d59f07625edda8df0c9d3d6, 168'h00f7027c029407ca619267eefd65408419add7d8a5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{258, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h009a984d1c7e1067811db09ac0e432b50bdfdfcd3b, 160'h44432ae69227c6262de5bb86fcb268ba58e0f805},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{259, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00a7a43e7ea768010355f0d8379a528a0e8109af93, 160'h7f536e774617d45674924d0e571b9c91665640e8},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{260, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h60123bd5b8bf38e6b9883fd8981f9e8189cf17a6, 168'h00faa772f9f27ad7a646bd95a189f59f1856a406e2},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{261, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h25952151a5fbe15c4184a0b1f212a8710f51d665, 160'h63c69705d2e525b5533bb545550d421f65a811fb},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{262, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00e76f11a18fdfcdb0d29fcec791cec461cd407348, 160'h35d35e84a7231179e3c90e2abcb463adfa0b2b9a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{263, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00f68c55d307bff3b43d41717624a9595f2d85c4ca, 168'h009f295ee2757b951b7c5b33cd9be3edc64427fbc8},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{264, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h779f3813ee80326bc082750b97ab9a32aded3451, 168'h00ffc66bac139a5cad892ff9df4e29476873daa7a6},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{265, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h5f1614bd3ed8ff1755186b3a16d0b46c98d4363a, 160'h70fed0fc130a3e15086d3dd5150b452cc9234dc2},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{266, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h7579791e611efa8183708f49f474db39e729201a, 160'h671ead3c5c8a57b90ce81cafea1cc7ac5c60018c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{267, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h68216e77a1c01777341e36782e4b350acf54fb56, 168'h008dac1469cf30f349f38b372ec879e989e1172aea},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{268, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00e3a395a24d5ccf2974fb2c07099f00aba3b673d1, 160'h437d95da3571611f9940c0ff1b3b29be5e65040e},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{269, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h0ecdf9992b5ebbee6770dad3aeefaceabc6106ee, 160'h5e849ff0607952682b51c8889d4b1dc0371f47fe},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{270, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h178bd60ae5c02fe00f058e4174535e62caf9ab3d, 160'h631242e73ef54d6e44a5adb7a1119e0467b52e50},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{271, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h755e6da6c7aebfec7169771d70aba265bbbd94b7, 160'h00c19262b7cb5e3be6a4128e54b8ef756f3c9085},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{272, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h7ec65c17c976fdab34e41858e39a48da52168e87, 160'h39df46e7912443837e38dbd210679ffc2be55d99},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{273, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h009b802f1318bf3fb0097629781da42684f0858660, 160'h0e83837218c15f2cd3a5c3ef9aab5e4b18f02a44},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{274, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00b8fe040f45392eccb25c4e8476928d3c2279a0a8, 168'h0098e144a6519e63e5772b707903aa9882865ee8c5},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{275, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h46591cc99953bc95bd791df1d49852ff4d155933, 160'h719ff20f870dc699c20be7add0701c6ef9f47c28},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{276, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h009aa5d6010f490139aed60d538e31381efe817d28, 160'h412d4d6188532313f22fc7a74ae9bf03f394ec9a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{277, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h2fa46053a3f59aefc91b4b286a15c31205812bfb, 168'h008453d2fadaacdd7ed6f7b7623915cc96a410f46a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{278, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h42c1dbc859090702b337f06304c32855aa032d58, 160'h54eb0ee6de7a6a75dbb3162a320d02433706fe5a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{279, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h7e868c5db1d0888024a6b360f4f911321a24e1bf, 168'h009e7565e15885b2962486d5c8d55669175d55bc23},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{280, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h6e4fbcfa8f008eaef72bf80224575cf6e0d5a6c3, 160'h1ebe3f075dee784663ec14b687aa54384078b8ae},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{281, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00aa7cecbc8ca25699e9ea4b84eb6868f21fec3a78, 168'h00bec86ae3ec814ca8e3f74a9db49c7800e096f012},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{282, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h72526c3ead0bcdf74e527c5498cf1b1df7d8524e, 160'h0b297ed48051140ca2ae592da02dd03e5f25ad84},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{283, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h46d3288ff12675c344e71be290d4e2d765500f02, 168'h00f7fe700a0c4758da1252a7aded14f61aa798694f},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{284, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00f1fc30dad8c322138e43d5f2b7555a7b34639523, 160'h66857f71e977375dde180754c15bd40b86f27eae},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{285, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h758a02aa0f79ff94b7b56086f803688072aa25a8, 160'h281a5a69e4571646333cedb80ed565d11a30f964},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{286, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h2660d3799b942b3e300bf7197f79724ddcb1ce47, 160'h3759b27452ff2465a0a947a904d3812e31405362},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{287, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h68279be7512023116b41e80143099f587731d960, 168'h00ed01510c3cc2db951c3b7e4f54bb0728a60219f6},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{288, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00f141f6fe5e020e4c01bbdd78dc326fa0d2c8860b, 160'h372afdf1cf524eaeeb62f195da1aef56c9c278a0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{289, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h0091161ec51b94f7adc6499675c4b508a69cde2728, 160'h41f90976b1dfc4e7d59df541e7e43904f3f0404e},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{290, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00ecafaa4a37764b6e3119bd06b44f963fd4db3bb5, 160'h6130126a72e1057006c865b626b91790fc90e537},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{291, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h008d72db18a44fa66006f2324d66ab8a86fc28a24b, 168'h00d5286dc61d445beea7952d30bf1f32ff725be47d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{292, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00ade33a64ea8e9dd1badd0e203f0f13e3cb3d171d, 160'h23dec9f58ab8f001126523ed89b1a7fb494c5677},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{293, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00ff4ba7ba455552e64eb56dc8872d10fed09a61da, 168'h00fbce266e3f340457d32650cf8692f88a74cacaa0},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{294, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 160'h2d7b0652f46d1cbe8f4a4f7556cb2d97f419d722, 168'h00e0a5718e218efbb22087cea30de8a4daf01a9969},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{295, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e4d9ffe5ec17db4997519d0ae4219c47d8104498, 168'h00b1ac39296f239bb18008b6711545873c9fade258, 168'h00843979d21099bda2c9f77bcb3fa8afe1f8a623c7, 160'h052a099c3aab4281b854ea672d22b3129de15faf},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{296, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e7e3adecd744fd9287a3ea9db7aef433855eb947, 168'h00c15fa9e3b893f09f46c54b4d20ef0ecd2666877e, 168'h00fffffffffffffffffffffffffffffffeffffac70, 168'h0100000000000000000000351ee786a818f3a1a168},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00fa19aff61dccb4982a520c4a844210d88245e643, 168'h00cad5c9f87432f65dc9609b50ae80da751a86bd32, 80'h351ee786a819f3a1f4f5, 80'h351ee786a819f3a1f4f4},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=80b(10B), s=80b(10B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d96a3a9da3eb41885ef8e6c1e1d59bc658c483cd, 168'h0088684298412c5eeaa9c8b20d15d0dc25d232b768, 40'h010000538b, 168'h00b95a110c2891cd3eb34a61499b56bdaa10ddcc4c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=168b(21B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h0dd2d6ce794df00949356bda4ce5933b41ebe45b, 160'h71a799413369c351373f18f66ee5ec3f08986c91, 40'h010000538b, 160'h46b6470dc8b43a7f5fe139ec959eafa683f28f2e},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h74151122fd301dec9139e1277de1063810fcf9c6, 168'h00f1797e4233303f7279e8bff017466a2963da7b53, 8'h03, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00af1ee8e681b5db8479ad6d2c3cce1bb6da8c87c3, 160'h427c7f8dc4de05c78a0ffcf5412ef343bb137e12, 8'h03, 8'h03},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{302, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00bebde6a1518a38bcb7fecfb6e70d92ec5de9e2fc, 168'h00931816f21cd2ff7c7317aeccf50a994a6fb44c71, 8'h03, 8'h04},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00bebde6a1518a38bcb7fecfb6e70d92ec5de9e2fc, 168'h00931816f21cd2ff7c7317aeccf50a994a6fb44c71, 168'h0100000000000000000000351ee786a818f3a1a16e, 8'h04},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{304, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2491a770160ee0f5c4964e3e361015b325e7b55c, 168'h00afc2886ff00714e00a1e002c6541141ceffba2d1, 8'h03, 168'h0100000000000000000000351ee786a818f3b477f2},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c7a2767e0ee2fcfcfb9f5956728977d6cb976a37, 160'h11627527eede9dad36f80302c1d39e5707674107, 16'h0100, 160'h4e9d3a74e9d3a74e9d3a8539de479664630141b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=16b(2B), s=160b(20B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h32c14d92c5bbf6e3440c4428bece01c77c4c847c, 160'h3cf05f2e5c56e67c8e583d982b6b4ef498c1cfdb, 56'h2d9b4d347952cc, 160'h6b725fdd61cad3a932f93b73e8fb939d7b7f98a0},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=56b(7B), s=160b(20B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h7115629c4cec6ecf0a96480a8e31326caea56804, 160'h2c713ebaaed6f69a15ef1eb5a79f38be468104b7, 104'h1033e67e37b32b445580bf4efc, 168'h00da25da25da25da25da26076a060a27a5b2b88c8a},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=104b(13B), s=168b(21B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a9309d2aa0520e82039cac944ec6ecdf2f830889, 160'h4291efe0efaf29d95e041b1a423a3b4f4d30c507, 16'h0100, 160'h3cc5990d6ad0679254b205b6210dc1204c382e92},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=16b(2B), s=160b(20B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d500ef5c55e6df67dcd941dad4e138ecb5ff7455, 160'h7d239fc8d9d3da2b799ed6c51f2f542f650eaecc, 104'h062522bbd3ecbe7c39e93e7c24, 160'h3cc5990d6ad0679254b205b6210dc1204c382e92},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=104b(13B), s=160b(20B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c2ac99d7f5028c94f65136175341d5366c3bcb17, 160'h332ab40a0de752e9c9509138f37ebc5761776977, 80'h351ee786a819f3a1f47a, 168'h00aaaaaaaaaaaaaaaaaaaace149a59c565f7c11647},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=80b(10B), s=168b(21B)
  '{311, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2805fbf5352896e2fa4d0ce04a1e46a1e0a54958, 160'h7d14fdd85792bce2592ec6e3adfab1232a1e1eeb, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2805fbf5352896e2fa4d0ce04a1e46a1e0a54958, 160'h7d14fdd85792bce2592ec6e3adfab1232a1e1eeb, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{313, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a02a7443fdd15c807ef45ce97a35b11d1d0ebcb7, 168'h00b224b97f6ddaf528d5772c0e27642c44ec79ca82, 168'h00800000000000000000001a8f73c3540c79d0d0b5, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c6613369fe141def6496756c4cb5235ce2dc043a, 160'h31f4cbc9d02e54433fa0772bae26cbd23779bb1e, 168'h00800000000000000000001a8f73c3540c79d0d0b7, 168'h00800000000000000000001a8f73c3540c79d0d0b5},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{315, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h76ea9df5b297e619a49f8f0286fa8aae73ecce6b, 160'h040250cd1f977f1c6790eac49704e9a3a3c58202, 168'h00800000000000000000001a8f73c3540c79d0d0b7, 168'h00800000000000000000001a8f73c3540c79d0d0b6},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{316, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h72d6561a598603b7b9313156aac55b41aa825cc7, 168'h00f340ee7492bb884bab5791726e7fba478e382819, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6d697574a79151bc53ba024c16b37fe6b87778f6, 168'h00850271deeb76262831378228ec4275aef3e21433, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 168'h00894b5a17a0c6db3c2579a652a6c80c6be6d57350},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h300cc0a40c609362f3f20b7c8e57a8f99e592436, 168'h0092a393c1bd3cd2792ca45b8bd56e4f7186817a54, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3b77acea21da4d7940fe4c7dc0f3efe476f36dfb, 168'h00fbc51dc5b9db0ba7eeb759786935cde5cf4b0618, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 168'h00aaaaaaaaaaaaaaaaaaaace149a59c565f7c11648},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{320, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00dcfc949a2a2bd5a39a8f48b0de700ab08dd59392, 160'h756a23dd5ea2ef12145c003267284a5b675a0826, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h7ce6e1f81fbdb6ebf382414e62c1c14200249a82},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{321, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c36bf5f8cf813744db69caf227e8c224eb06ca03, 168'h00fb4187818249d1b14c1485d8d3b4c8756138c89b, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h4ab240469b50549275e2e01f81c8728b51a53628},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{322, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h355ddd7796c24783c9b55264be1156ef5f76c568, 160'h333126d0e19d66868545c91b193a33018395a678, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00a14d77e73be9d42f3f4eec1e2aec1f4988327bad},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{323, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2df2324222c2a34e1988aa4cea44225d5137ae9d, 160'h5c0033b715b1614b9375f7addf8c2d0a2c1b9fb8, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h57dc8cdfdfb0e210894b6c52e53ff10907c71962},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{324, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00ce705444a03779bfcdef89d67ec096098ed63cea, 168'h00c5d9a58ce038b2fbc5ec13368a40590d39c1ade1, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00c8cdfdfb0e210894b5a1a3b75107ff8b538337c1},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{325, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h11e3b7937ae51b7a419529cf955ce7de33c38f20, 168'h0082d16eb3f27ab2f880884d93dfd09d6f300da51d, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00919bfbf61c4211296b43124fba8956fdb364ce17},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{326, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00894a29444a70a0eb5ed46a353512fd2207048b0c, 168'h00f8e70a6fb6cb6816c007d00c286e43c3f590212f, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00dfb0e210894b5a17a0c709a6c54fb9a74cf9dfcb},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{327, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6ac3a901506eefc03beea1c282cb6696326e48db, 168'h00c9604ed9ba2282eff1412f37806c10ecffe8aefe, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00895d39009004bc13b7bff51e58acd24066a2e37d},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{328, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e44f04c7f8a83e3acfe938434bfffe8fe73663ef, 168'h00cc258bd2d073b7a9c28b791887476eae2e249e58, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00da8789025ce0af8603bf87edc9e62151f396a644},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{329, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h705b3a456cb6e36cf5dbee426e0665b12f35452c, 160'h3e21f76bba44e797f86ee316080b028979163935, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h0083191e07e04249140c7df3d084c4e6d6f37d06e9},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{330, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h1602e1a8185f83a842ef7eac0fa72c11a1033a92, 168'h008930f9bacd398f87462be0dbe38c6dc36426a8b1, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h44a5ad0bd0636d9e12bcd32953640635f36ab9a8},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{331, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h5b52a108c602cb117befbefcaef469b0a393258c, 168'h00a15232d2a7d22160f217b7caf1410b66d9978abd, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00d0a6bbf39df4ea179fa7909e893963b13dea0e8c},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{332, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h40ff772b7e38ccfd01bc7ba94938890e1ce09678, 168'h00957ff3dd0c66ffd5f20c1979ab8ef74285c544e0, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00aaaaaaaaaaaaaaaaaaaabc5fa28238085135e078},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{333, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4c4160c33fd9bb567628218d0233dc8a9b220b63, 160'h4d8fb88de219a3f539a0eed7a25f83e3a339c08d, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h6b4aaa62e57733898782c2fc5c2786bed659b644},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{334, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0086057b5f1c0ac3682f375517184d9d098e97c870, 160'h532d07fce6031da8c92385279a8d45955c07b731, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h58f915945cb8f92c33b91a69f8efb78fea695455},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{335, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h68db60c95140e3fd8eebce400a806622122b1ce7, 168'h00887c0655a0c3af94b128be056561444a96c1d366, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h5630164b8c5d7636000011e25c32facb98cac6fc},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{336, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h7a9effc019cb530aa9225231dbbc25545817e06c, 168'h00da9e301fddc37794f989549bf63508a731d50754, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h0164b8c5d76360000000004a05513b244cc73c9f},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{337, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e9666ddd4f967bbe098f6b8e4ee43152241f0f44, 168'h00a906666bdaafc897e7a145aeb6f08ea88ad119a6, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h02c9718baec6c000000000940aa27648998e793e},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{338, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e547664d205f9fff721e515031b2cc2b3c91cf16, 160'h6b068a123ae01160608040675422ace4462ff99e, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h008c5d76360000000000001d204b5f683485b683a7},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{339, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2d5284de38eb2fe49a5a2f972ec865015f50d64c, 160'h54db02f299315f526b5a3a6c1dc7a7f4cf3fcd1d, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h618618618618618618619b98b30bd6533e0a9093},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{340, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h5c270156584fb1d0f7aacafe3b8610a95de3ce5a, 168'h008c25025900de5354f04aae6b77d253f659b1770a, 168'h00fffffffffffffffffffffffffffffffffffffffd, 80'h054fe3f3dd9c185cf68b},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=80b(10B)
  '{341, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h33bfdad102d60c52addce3802abccbc7dc3c7956, 168'h00db4ab15fc608ff386121022bcf2c3ea06d387b42, 168'h00fffffffffffffffffffffffffffffffffffffffd, 160'h5555555555555555555578bf45047010a26bc0f3},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{342, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h0a01ffc9638f8734559ab2371dc4b431a9238304, 160'h0925e3be4f7e5007b2ced6e6dac3a9cac02c566a, 168'h00fffffffffffffffffffffffffffffffffffffffd, 80'h1a8f73c3540c79d0d0b7},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=80b(10B)
  '{343, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e0c407cd8d8b3507e36c0aa8e15b4f17f9e07d72, 160'h667946f46d6c618b628c048b3fc808b2c40e31a3, 168'h00fffffffffffffffffffffffffffffffffffffffd, 168'h00ac7c8aca2e5c7c9619dca7c4703b2fd46f057ae0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{344, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h74d02bbd2218bb4ea9492df5ab596cdc77d81f96, 168'h00bdd4a5d816ab10076b6694492608b85851704a30, 168'h00e278b476b12f0dfe75e1616063ab70f40e7a7b2f, 160'h71c197e44b684b3b8f972367caed38b40c9ee4cb},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{345, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h74d02bbd2218bb4ea9492df5ab596cdc77d81f96, 160'h422b5a27e954eff894996bb6d9f747a6ae8f6243, 168'h00e278b476b12f0dfe75e1616063ab70f40e7a7b2f, 160'h71c197e44b684b3b8f972367caed38b40c9ee4cb},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{346, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b126e61fb24c9932a12c50a14844887677276bca, 168'h00d4710b84ef34a8b28e290179e864ab350c761785, 8'h01, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=160b(20B)
  '{347, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00871b534b25d5738f44c1943c8b634ccb7444f1d1, 168'h00b581ccae151d819301047f0442cbb6756b40f82c, 168'h020000000000000000000000000000000000000000, 160'h333333333333333333333dd2fb1aee6b63ed2048},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{348, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e0c8238a5ab89f192a0190821b958986103d0966, 168'h00bd64baf7e2417212d99b4a899264e122db67e99b, 160'h55555555555555555555670a4d2ce2b2fbe08b23, 160'h333333333333333333333dd2fb1aee6b63ed2048},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00ad4577f7f3008aa5ebbe149509ad3de4b7bac270, 168'h009f1a6ba48149bde27ebf3a8fab4b8483676b4c95, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b96c963f6c4c8677f0da769772df576c56876b0b, 168'h00fd93bc9cf6f640e36342c764ad9ce5e8fa86c3e3, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 168'h0092492492492492492492677f5fbaa932d45c5c3d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h008779d9d40470df9c4b6c53c27330a0f0c748c01f, 168'h00abe5c16182899fe3d702ee89bb14a51aa8ff6cc7, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h666666666666666666667ba5f635dcd6c7da4091},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h0d70d01018f55e36464782339c2c8f4a1b963738, 160'h34d124028d77ee31fe2a3e2c10c2a4f7a5fa0dde, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 168'h0099999999999999999999b978f150cb422bc760da},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a7afd930bd9f9392483245ccd628be428e0f6555, 160'h36c945fee505c5fe855187ee725402995cb0e701, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h6db6db6db6db6db6db6dcd9f87cbfee61f45452e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h45fb936471ddf35059c571f794b7fd6f23f752ff, 160'h3fa9603f8c5a370da68f3f812802f0da5d21af74, 160'h26788d2ba41a035954dd638d883e136ab900c8cd, 160'h0eb0f1bc9eaf6ad85b2d94e5e1b53937df61a288},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h49d0064ca551c15fac3f13f9cc44a8309c31e721, 160'h3d403f3bee9ceaa243e492cb9a8f83e92c3c11b6, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h55555555555555555555670a4d2ce2b2fbe08b23},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b08fda3bb59b426e374c3ed3a7eec174379904ad, 160'h72feb9fc39221407859eb30c1a1166aaabcf5c15, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 168'h0092492492492492492492677f5fbaa932d45c5c3d},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h491a910b75f57a4cfc2fa7c878c0a23a725952d5, 168'h00aeeb19e0aba884da4cd64574e785ab9323d0f681, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h666666666666666666667ba5f635dcd6c7da4091},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d7f1c5d7a03ed20e786e856e666184f2ca541aac, 168'h009eec69b468ecb87fab4cade385d2bd9fd762308f, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 168'h0099999999999999999999b978f150cb422bc760da},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0099704a8b543c9ee06a913b9476d6e1b741e28368, 168'h00df8cb71743ef9903231dcfeadcacb4e640192397, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h6db6db6db6db6db6db6dcd9f87cbfee61f45452e},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3a81a3afa818e6511baed5c8d52c617223cd3608, 168'h00f3f13a8c30bff4cbfbad5d0789f8e12bce995b43, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h0eb0f1bc9eaf6ad85b2d94e5e1b53937df61a288},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{361, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 168'h00feaffef2e331f296e071fa0df9982cfea7d43f2e, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86, 160'h2492492492492492492499dfd7eeaa4cb517170f},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{362, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 168'h00feaffef2e331f296e071fa0df9982cfea7d43f2e, 168'h00894b5a17a0c6db3c2579a652a6c80c6be6d57350, 160'h2492492492492492492499dfd7eeaa4cb517170f},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{363, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h0150010d1cce0d691f8e05f20667d300582b6d45, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86, 160'h2492492492492492492499dfd7eeaa4cb517170f},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{364, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h52dcb034293a117e1f4ff11b30f7199d3144ce6d, 160'h0150010d1cce0d691f8e05f20667d300582b6d45, 168'h00894b5a17a0c6db3c2579a652a6c80c6be6d57350, 160'h2492492492492492492499dfd7eeaa4cb517170f},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{365, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 160'h46f1a7493b131f3c6032e9612b8e1bd3d1a3104c, 168'h00e3cef3c8020c277ba45bc93a9a364f07eba8302c, 160'h2b5ebaf4211158c687625922bd903253892cf834, 168'h00aed36914690e0d99637b92439539a13bd8e6d800},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{366, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 160'h46f1a7493b131f3c6032e9612b8e1bd3d1a3104c, 168'h00e3cef3c8020c277ba45bc93a9a364f07eba8302c, 160'h6d8624bff7719b53dab811bdc0e434a5e9f02e8d, 160'h0b50e6dce0f5c1a757290eed8df0aa8092b2ff90},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{367, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h46f1a7493b131f3c6032e9612b8e1bd3d1a3104c, 168'h00e3cef3c8020c277ba45bc93a9a364f07eba8302c, 160'h2039f168a3a1f9f0a3ed4f11be9d5d0a9807eb8c, 168'h00ca18c2ebd6bff0ce46dcdefd16ab455fb36391d2},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{368, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 160'h46f1a7493b131f3c6032e9612b8e1bd3d1a3104c, 168'h00e3cef3c8020c277ba45bc93a9a364f07eba8302c, 160'h4f71a123bf7c4983f5707c17ce4782c833e833f0, 168'h00dcfb123cf5470f21375e62ba4054ffd9a836908c}  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
};
`endif
