`ifndef WYCHERPROOF_SECP160K1_SHA256_SV
`define WYCHERPROOF_SECP160K1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp160k1_sha256;

localparam int TEST_VECTORS_SECP160K1_SHA256_NUM = 227;

ecdsa_vector_secp160k1_sha256 test_vectors_secp160k1_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'h00e0348c201105978ee3ab9c565cf9a63261a58173},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'ha89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{3, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{96, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 184'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df230000, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=184b(23B), s=160b(20B)
  '{97, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 176'h1fcb73dfeefa68711c561ca3b9e60568687135400000},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=176b(22B)
  '{101, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 184'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df230500, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=184b(23B), s=160b(20B)
  '{102, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 176'h1fcb73dfeefa68711c561ca3b9e60568687135400500},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=176b(22B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 0, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=0b(0B), s=160b(20B)
  '{118, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=0b(0B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h02a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1dcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154dfa3, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1fcb73dfeefa68711c561ca3b9e60568687135c0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 152'h1fcb73dfeefa68711c561ca3b9e60568687135},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=152b(19B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 152'hcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=152b(19B)
  '{128, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 32944'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df230000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=32944b(4118B), s=160b(20B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 176'hff00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=176b(22B), s=160b(20B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'hff1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=160b(20B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 32936'h1fcb73dfeefa68711c561ca3b9e60568687135400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=32936b(4117B)
  '{136, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h01a89cf5aa14f3e5d8a031291bddafd4b93b6b95d6, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'ha89cf5aa14f3e5d8a02db727aff07d83a73e2870, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{138, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'hff57630a55eb0c1a275fd08fde392fd6e18eab20dd, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h57630a55eb0c1a275fd248d8500f827c58c1d790, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{140, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'hfe57630a55eb0c1a275fced6e422502b46c4946a2a, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{141, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'hfea89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{142, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0157630a55eb0c1a275fd08fde392fd6e18eab20dd, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{143, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'h011fcb73dfeefa68711c57d59dd0c5b1033287ebf3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'hff1fcb73dfeefa68711c5463a9a30659cd9e5a7e8d},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'he0348c201105978ee3a9e35c4619fa97978ecac0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'hfee0348c201105978ee3a82a622f3a4efccd78140d},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'h021fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'hfe1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 168'h01e0348c201105978ee3a9e35c4619fa97978ecac0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{153, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{157, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{163, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{167, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{176, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{177, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=168b(21B)
  '{180, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{182, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{183, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{184, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{187, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b3, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{190, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{192, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{193, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{194, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{195, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{196, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{197, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{200, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{201, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{202, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{203, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{204, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{205, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{206, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{207, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0100000000000000000001b8fa16dfab9aca16b6b4, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{210, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{211, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{212, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{213, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{214, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{215, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{216, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{217, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac73, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{220, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{221, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{222, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=8b(1B)
  '{223, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h0100000000000000000001b8fa16dfab9aca16b6b3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{224, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h0100000000000000000001b8fa16dfab9aca16b6b2},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{225, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h0100000000000000000001b8fa16dfab9aca16b6b4},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{226, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h00fffffffffffffffffffffffffffffffeffffac73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{227, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fffffffffffffffffffffffffffffffeffffac74, 168'h00fffffffffffffffffffffffffffffffeffffac74},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{239, 1'b1, 256'h9338b2ec2eeef8c37432cdf94086f4e6988a80db24816c0d4ebd0175cdf55632, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0097f6ec6b77f27688037564fb65fa69190a4e8d4d, 160'h10f26104009337dfdc87787c430052985758391a},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{240, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h19028f9da4be925a155ff4fd71ce09058d3ddfcf, 168'h00fd0c0937f65e6a8b0748c785d1ccdd1c2fff2759},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{241, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h2e63b73510882b93c69a8d00767f9b9897262b2d, 160'h2e401df2d03607e9a26e16f9550abbc4d40e888c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{242, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h4296974dca1d2ac6db892b65e2ae5877ab243e1f, 160'h35b0559258b7be92dfa2575d78c9798058e16a4e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{243, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a4503b37879fc1c8c49fa1cf0fa66a6eb2ae01f9, 160'h636d8b378af14b81ad610f82f6ebabdca927bde1},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{244, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h0766ca1cad1e6e47a3dc8d86d8ccc18624498273, 160'h47791918c5bb5511cf25194fd52d7cca97a931b5},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{245, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h71637fa756fcbc3b8313501c1e651569733ee71a, 160'h12334122b218782a145446996546bcca95c7c968},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{246, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00b7969db89f2ae5fda32dd732d604c44a5978c368, 168'h0082fa4d1c095cd8ca0fac77f6c9bd554f2e498b0b},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{247, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a1541f7355f7d2f4cf303874ae692be3dc1ee772, 168'h0094c4b5f00de0d1917f465c1e46398160adc2569c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{248, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00b1b688b3d205d80decb43976513a5bcba623fd6b, 168'h00f6354d422014c47c2f917ef2e2e12f3dc5a74156},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{249, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h332bdb558a26d7c8d157c2ee72052b1e759b2739, 168'h00ebb2a43926bcb47e57ccaad24411ba6e9e08a474},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{250, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h6cbe031b8dfd5142eb7c8f69c9d4d3f25f48a903, 160'h27685c54fd837ac971f198b661620eac851d9d7a},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{251, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h009a91b10985e3d766c7115a63fa166166302f3ee6, 160'h7b6f264c4f7e47f16d966377417c4f7edaaac6cf},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{252, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h008a84181b7ed1a6092f1df4f8eb9b9622a802db5f, 168'h008b5f4e66ed1a8710eda97f37d452d3384d5fb864},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{253, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00f669f4374b1f9aeec9a38469653019721f76135d, 160'h24632ae6b502d87d185a3f78d1ee4c94344f309b},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{254, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00edfadda70d827712cb8f22383892a04878dd25df, 168'h00eae0caa9985f8bf391613637a7ad6bb295ecd7ee},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{255, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h008695d692e98dc81f765a287733b5947da8769fc4, 160'h5485ac28d4694fbcce00b362846489b8aee94104},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{256, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h5b58249bb9fc858db67257a4bb5d21df6d8a1dc5, 160'h74d16dbf41fd4d5bd148a0cc020f6ea6bed1d5eb},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{257, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h46fa4b37d994ede647aa00e8552867a0fd932c25, 160'h75a0850d1e7d0d0e3a796a1df069d5bb9eec7309},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{258, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00ae613edca490cfba96a489081b3f539d89058655, 168'h00c393f881019c5b7612e48c1e44ecb10847605e8c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{259, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h008bb6449c147d6132193bd7f9a6f33573083dbff9, 160'h7a0c45cc495c000576b4bddd059db28408e52d59},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{260, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00b4b1920e46371d08090a28f2a8ff1a2f909acd5a, 160'h590e62faa9a50e20b308cec56b686196ad95db96},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{261, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h009725e0058731608d09d96bcb3acf8d8b802cf396, 168'h008d360949c7ae08b6536fb6904f3a5c922e32a216},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{262, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h514b2af7da92ce789e3eeed98044699530e5af30, 168'h00e606484cb7d347843c64cff2518319108e661094},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{263, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h6e3f020af00d2b56ec3e92b23e981486b679bd44, 168'h00ba5d05d594bdf5f84fc1303963836fc09538c7ba},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{264, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h30894ccb595c048cb6ff9dcc5b974b5a72e9fb95, 160'h1c3b805772e98845dbc660d3675174e9842c7f2b},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{265, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h6de326ca60d74a5997d4137b4b6f66f9a6ebff91, 160'h6a5f5b88569920c4f7644a476280a6e711ddf058},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{266, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h4322df2ee1b393f924d41087fc8e1192a78d4d81, 168'h00e1fcb8341b8746f6e286344c4a6568fd2c29c478},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{267, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h5549776bb880140a441ac4d694bd91c683b2963e, 168'h00c0238343c8e2cd3938d3a0c9323ca4e900a60e0f},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{268, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0093b97e687275cb1f25f21244b0deb68a764e670c, 168'h00f273675cb6c96cce93b58b83276bac609daff217},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{269, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00f7e0342fd8e29e0b750d494b0196989692bddb4b, 160'h7d161fad96dadbbbcccdb20c9f824d58989570b1},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{270, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00eaf1f3c050520411276b0be225a15d3986bbf065, 168'h00c1c393f5b9f1e2c554bd4669da940b8a27b33d73},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{271, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00fcb46239790add12b1a45bdf6bbb6a40dc552b1d, 168'h00a4fe379b92ce6e25e5d5ff464b1adba0113a63e6},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{272, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h39f9b38cd943bcc3ca0d47a276c419e1ae94643e, 160'h59027aff40966014bdf62c7f6ff1197e5093644c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{273, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00f0aab4b3d38ed8319769cbd68fddd42801950d5b, 160'h1d83776d13eff23faa7186f4f24e866f0ba898d8},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{274, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h193ee899b803a67b1828a1ffc0f10e1c6c107732, 168'h00b126655e5416b012d7e79abedb8c8efc0e77cac3},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{275, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00aa38d9765ab14baee6382e3a42dcb1d0070ea37b, 168'h00989d56b71e597146e36226851ad91fa8535dc1f1},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{276, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0085d763ddb93a69a1ba30a32d8f16fdd23be1922f, 168'h00e74a2f24010e0d608447226a3095b7002a60c79a},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{277, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h21b3076b15ec039137a36b158f4b6a14cb6c340f, 168'h00aa819af1d2df1592f5ca4e2a0133d2c15018df1b},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{278, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00b9ddff30cdc294a62e3b7135bf2acac7f8afeb95, 168'h00b9757d6f4f181702bb43ee6295bec560db7f941f},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{279, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00b45fc55b99384e7e929aa43d017e398b61ecd034, 168'h00bae8572ad844856b0827e201045ed8580af05806},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{280, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h319a4b68b6e8b6f8ae809a690741f11fea657a53, 168'h00bd931f12b8f8853a8f7de98be48aa813a18ea3e5},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{281, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h0c09432e6d3ea9798dbd0d7411816a526d08fc1e, 168'h00dd1640db6439f6c56637abd9979b8652ea04f36e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{282, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h0083dc9d0bc5536e759195551c29e8b3343c069499, 160'h0db4e57490659d25c3202cf9c525f8dde99466f0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{283, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h640505fe143986f7b46b80ec44d83c7b048a34f8, 168'h00bfff5d4d604a08ffde84f518998145a277ec1376},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{284, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h1c77e9430c235c33a93d7f74ae2b1b67afb75191, 160'h4b1b6c4c49ad002a1017e5017fc495a4ecc85c1e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{285, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h2d3a0bba220b15814b0cac3f1a344f648755ff8e, 160'h68f067f05edd4b543a0d8a92f5a6025769617029},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{286, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h7008b9ad8a2d21857773a74eb2646c5f182fa972, 168'h00e093cd77398b29c5f40df9d3b13e9a84f2e92c43},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{287, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h3174c392114a6e623a4778bbd26dcb8ffd0a5e06, 160'h3425b221031c23d6a99efa813109e53fe5402176},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{288, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h009b2e4e552cdebbbc0123dd165d199a77c1c36328, 160'h3f8395fd386efe25c512708d3536d5559604e41f},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{289, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00c1f62927ac353ddde5a6f95244aac6dcab007ef0, 160'h70190e74000a2e8d23321d2c2cdaf640b3831923},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{290, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h16771ee4085694c00ee10b616484d87e878554d8, 160'h67dffce5c711eca8e370d2bdce36aa0205e7d313},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{291, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00e742767507f2aba4c70b931201b3466a87e321e5, 168'h00948c505631602bc82ea74d886171a90d67364874},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{292, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h26177ce30103120b5d24eb052797e5b2b9d31f0e, 168'h00b8976208a7b7a27cce87abdd55924a9543138552},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{293, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 168'h00a78db1954f1ca4dc3766a6d1a14757610573b78d, 160'h36da520ccdaa9da29751948d54636e6474409327},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{294, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h62aca5e281c1fa6cdbb65ef92897c2ff5226b3bd, 168'h00d0b82f15239a0d7c4b04a6537dfedac69571663d},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{295, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h1b1fa19f5645059f46ec5aa9d033628f079f3218, 168'h00e2809349c90a70bb00304b52bf31ac028c3dcdaf, 168'h00fffffffffffffffffffffffffffffffeffffac72, 168'h0100000000000000000001b8fa16dfab9aca16b6b0},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{296, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e0cf91de379ee7b1a36dccdb7741b600e23f2220, 168'h00e035f7b0c969c775c8dcd93a41622ce1e37484e3, 168'h0100000000000000000001b8fa16dfab9aca16b6b2, 168'h0100000000000000000001b8fa16dfab9aca16b6b1},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=168b(21B)
  '{297, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h66fc1dee23644d9e110c2be47ae70679aa0dde2b, 160'h5d2db956ac41c8f82463ee013d64067d054516b9, 168'h00ffffffffffffffffffffffffffffffffffffffff, 168'h00952d47af4507c04008f3a63ff8f591054f3dc5d5},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{298, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h147bdd2b325d3a1a5819585c5863478144ca08c6, 168'h008523348abbfbe3596a2e182459f699b9a86c8c42, 168'h00ffffffffffffffffffffffffffffffffffffffff, 160'h6d534720d85cd391e0a69b6f97d70d4df0b01bcf},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h012a78f3ceb2c5606f824b90b4151a7cd788c3c8, 160'h6216521c8b038e7080bb5601ac8b49e96826368b, 8'h03, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00cee7f5abdb03bb603a30a7a781d2249708931e28, 168'h00f459dfe37fef1cc13d5832452381cc179e708728, 8'h03, 8'h03},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h48c7400e22d2ef7354b820eb662105e1b6e44a60, 168'h00a329f8bd69afd5aa91d4e18d3cfa2428930dee68, 8'h03, 8'h04},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{302, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h48c7400e22d2ef7354b820eb662105e1b6e44a60, 168'h00a329f8bd69afd5aa91d4e18d3cfa2428930dee68, 168'h0100000000000000000001b8fa16dfab9aca16b6b6, 8'h04},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b20b8d8201c0b40c80085361307f77715c519054, 168'h00dba52dab76d7a79bd4c129dcc945417dc1f03dd7, 8'h03, 168'h0100000000000000000001b8fa16dfab9aca298d3a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=168b(21B)
  '{304, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4e93629502fc5f1e2968ee25556e14f1d6fac057, 160'h7b892be36a100c193a9bd21f6542611a8c8972f9, 16'h0100, 168'h00bf7efdfbf7efdfbf7eff45d547891383e9d07c92},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=16b(2B), s=168b(21B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h079fdc2ba58d2ce63611b3459035261405e179db, 168'h00dc027bf8924259b02fc4aa144b7dcb58e60eb365, 56'h2d9b4d347952cc, 160'h415936395bb46f9943914f2100607aec6cf33d9d},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=56b(7B), s=160b(20B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00990cfd22fb6aacfd6cf03761c7e57aa2a5d777d8, 160'h5fce9841ca3a588d3a475e079971814d3ae9fa44, 104'h1033e67e37b32b445580bf4efb, 160'h6b946b946b946b946b9524e49d0953123b068e85},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=104b(13B), s=160b(20B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00ab206289a1885cc739095c9a40edd81e8d5b70e6, 168'h00b8fcf0d4a8ab3a5bfb2e0fba0a093a1c16339ebe, 16'h0100, 168'h00c9dcec4e3faba91b1d9b7af283de683c91475c19},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=16b(2B), s=168b(21B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e76b9acb3c2fe6f5f4846353ed5070886b25c683, 160'h6998969342fa39157ba598d281d3be12b987a034, 104'h062522bbd3ecbe7c39e93e7c26, 168'h00c9dcec4e3faba91b1d9b7af283de683c91475c19},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=104b(13B), s=168b(21B)
  '{309, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c0f30e6dd1e373525383642bd45c9c3afa50def9, 168'h00dc9d63fa05fd685623d5f3690f3de32335e6ebb7, 168'h0100000000000000000001b8fa16dfab9aca16b633, 160'h55555555555555555555e8535cf5393398b23ce6},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6b54692483b37d1cb63c0ba6b5c74af4fbb5b336, 160'h67ea2957b75513d2ae6d1a2ea9ece586da947c9b, 160'h55555555555555555555e8535cf5393398b23ce7, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{311, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6b54692483b37d1cb63c0ba6b5c74af4fbb5b336, 160'h67ea2957b75513d2ae6d1a2ea9ece586da947c9b, 160'h55555555555555555555e8535cf5393398b23ce7, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h38cbefd21b9c1fb5936dff37a1a56e69eab4aea1, 160'h75620f851c610de6566ebacff24799b292f062af, 168'h0080000000000000000000dc7d0b6fd5cd650b5b59, 160'h55555555555555555555e8535cf5393398b23ce6},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{313, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00ebe4094ffa91819212f388679a03cf71bb4804bb, 160'h2e3d3984d88b7a8672c5bc17bddbc6e6b6083975, 168'h0080000000000000000000dc7d0b6fd5cd650b5b61, 168'h0080000000000000000000dc7d0b6fd5cd650b5b59},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h406655dacc20bde5d98ad97aebe4c802b956d6ca, 160'h46414ac3bae4c1036dcf0be063499416c8a3b4b2, 168'h0080000000000000000000dc7d0b6fd5cd650b5b61, 168'h0080000000000000000000dc7d0b6fd5cd650b5b5a},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{315, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3f1ba8aeeae79f6d241fd8be46ffa6f3568723b1, 160'h1dc482a95568e8e6cf5025cbf5b8fef9ee4fba1b, 160'h55555555555555555555e8535cf5393398b23ce3, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h47a6a457ba4e369309e211e0ee107e52c5eefaa8, 160'h2236ef54f95d209f58b74adbf17cd416472c4516, 160'h55555555555555555555e8535cf5393398b23ce3, 168'h00894b5a17a0c6db3c257cae09057a136f93bf9de0},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h41f3d434600a3f8a8a31aebe2cddfe2bc2b0d6e3, 160'h133cd88bbc0a4d81603015f3dce1ea82e1fa49dd, 160'h55555555555555555555e8535cf5393398b23ce3, 160'h55555555555555555555e8535cf5393398b23ce3},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h534a6949f782f5d4eced5ba6631c12be9f379f17, 168'h0097cd5d75ef0cf2cef901a3dc4e1d9e033033ec4f, 160'h55555555555555555555e8535cf5393398b23ce3, 168'h00aaaaaaaaaaaaaaaaaaabd0a6b9ea7267316479d0},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c1ba77b68c24397599f5eebc6b4a48f4f8caf4c5, 160'h3786ae759de63750382753b333576f5c1b26c540, 40'h0100005383, 160'h7ce6e1f81fbdb6ebf382414e62c1c14200249a82},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h28a2173e9bcd94c46d5dd3d160c8d3c6f5f392cb, 160'h77ebe984b44814ef24d6d2570ecbea704bf587a0, 40'h0100005383, 160'h2e5c5c1b387dfb0e98740c28008998e351483cfe},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00fb75a1a2c846d22d787e73d1d7bc7c81b27ce6d4, 160'h4f5ca24aeedd2e6dc1ed2c55f59ef00ce44f800e, 40'h0100005383, 160'h34a4abe436ec3fc4d118f7aceec0df6fdae800d0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h04436adf3f58cab7a2f5dc07d207816dcb1ea7a5, 168'h00b3899f380ab7f9a8d385933ec57cac4291a7a6c6, 40'h0100005383, 168'h0086336155015c2560894c41430a3badaa67bd104d},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=40b(5B), s=168b(21B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b5594d926de21168b0f60962e720c7623563158e, 160'h47a500835967a864bcd75d14ae3780ca0f154895, 40'h0100005383, 160'h36155015c2560894b5a1d735e4fe734ef48690c7},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2df812587ffa67e82da47bce7b72446b7235ea74, 168'h009569210bcbb40d4fd9ce06d58f74b8ecc964bdfb, 40'h0100005383, 160'h6c2aa02b84ac11296b43ae6bc9fce69de90d218e},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e3011e8fb90bfdf17424d59d0f7c9757e0a9ba8c, 168'h00ab28c585258001594b87d83dea00294c4a4ee79e, 40'h0100005383, 160'h015c2560894b5a17a0c6dd93d9d5492d33928391},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c2fb0180784a8f5074304cb708002635e844b3d5, 168'h00c8eff920e00d4ba506c58ca250fcf641b18e6f61, 40'h0100005383, 160'h18f90d4fad917e9601713c4ea95ad2def7b0806f},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{327, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4b4e5f5747dbd6ff941b8e7dcedb35377375225a, 168'h00d2292389c374d7d22668c5b0bf439c585c11d649, 40'h0100005383, 168'h00da8789025ce0af8603c10bc8f93f24d3ca0bbb8c},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=40b(5B), s=168b(21B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d42fdd8bf04a07864f49cf7a63b1bfdd98f6de07, 160'h2f1de4511955122331be5c73e46969bc940c8d5a, 40'h0100005383, 168'h0083191e07e04249140c7f77abb41dea58c9f21c31},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=168b(21B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3943713524548260c840a4c833091e2682bac598, 160'h05acb1d6bca1c685ed1bca4d05dc6ecfb8f22206, 40'h0100005383, 160'h44a5ad0bd0636d9e12be570482bd09b7c9dfcef0},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4c21a2c434cac9188f48721e1d0b160d5e3d8502, 160'h73d7e1ccd671a4f7ad0b9b150d4c64a2982191a6, 40'h0100005383, 160'h1a5255f21b761fe2688c7bd677606fb7ed740068},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2d36e6f01f0646f272289d73500e4a2fb7450294, 160'h5500bc561c648880fe99476b80b19cc3dfa3169f, 40'h0100005383, 160'h55555555555555555555e8535cf53933ee07ae12},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{332, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h633842757a9dc3b198de959bc34cc10ac9539be2, 160'h14b55c72f731cbec1a6cc80c30c9a868dee85233, 40'h0100005383, 160'h49714251df3ec8f3a9f5a39c44e3be5e5fbfdec4},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h03688c836288d11d9978ac2cd41ed4884e074555, 160'h1d524a23c8b8871191dee13b6ed4b3dc8ba20105, 40'h0100005383, 160'h599e266b8075ef551833f964e68b1787c9a5d565},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{334, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h37bafb3cba163d05559ca3639906d764b3a213ba, 168'h00b30c713077a32dec18465e1e73568066bef58532, 40'h0100005383, 160'h77f11661e51ad7f10000ce9b8a9fa0b557fdb532},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{335, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c66d00b9cd6b5b5903b2ece209470e712b96f515, 168'h00c9748522a17b59a60e74c69d7de161a5f9ffb532, 40'h0100005383, 160'h11661e51ad7f100000001df88363f82efb0f9833},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00fe4479b039c9781af875e51a40a1988f99e4777b, 168'h00d4b01aa8430b9a6b271ed609cbe59ad97f189bf5, 40'h0100005383, 160'h22cc3ca35afe200000003bf106c7f05df61f3066},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{337, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h7a3723db1ff831198e0f78add2c3b1c3b888d444, 160'h125049ac5b9296d97a8989085f5e26f1b27a606b, 40'h0100005383, 168'h00e51ad7f10000000000018aa5f3d593de462e642d},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=168b(21B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h009d0ce306a8c0ae72ab613c6c300680b23a5093d1, 168'h008d096766e271f991f2d0d37f73b990480375ada7, 40'h0100005383, 168'h0093b13b13b13b13b13b14afa3f9810a631bf96631},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=168b(21B)
  '{339, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00db6a0bf3b46e770976988c7e90a9749c6921e387, 160'h6be8958d44945e9c7fff210906cde88d02674901, 40'h0100005383, 168'h0080000000000000000000dc7d0b6fd5cd4b71b966},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=168b(21B)
  '{340, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h142b1e76f507c710c779cd9ddbe7b26ce567203c, 168'h00f8face07dbd07b082d69b682443b9b15e15db739, 40'h0100005383, 168'h00aaaaaaaaaaaaaaaaaaabd0a6b9ea7266dc0f08a1},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=40b(5B), s=168b(21B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d09d259f08eef381512ece8c5022f1e368dae62b, 160'h31de3c17efbd3f13e8f8cac2546cfb6debf9ee3e, 40'h0100005383, 168'h0080000000000000000000dc7d0b6fd5cce50b3198},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=168b(21B)
  '{342, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c8faedf1be8ccfd14b2f1c140700282ef12ced9f, 168'h00c4a328ee1fd457cc71c14009225826571264d7d5, 40'h0100005383, 168'h00accf1335c03af7aa8c1ad92f7eb5619149de460c},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=168b(21B)
  '{343, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c49a2de709bf46809e0daecbc359de43e56728a9, 168'h00baa96a39b7f0fa137256ff479ac7d974e18bdd35, 168'h00a4b1717eddc1e47de4efbefed814f306e4da582f, 160'h1708da0962c5ea1895c30878d90f3e72fef7190d},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{344, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c49a2de709bf46809e0daecbc359de43e56728a9, 160'h455695c6480f05ec8da900b86538268a1e73cf3e, 168'h00a4b1717eddc1e47de4efbefed814f306e4da582f, 160'h1708da0962c5ea1895c30878d90f3e72fef7190d},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{345, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0098defbbf1a0a86d2cfee186065c697f65f471f99, 168'h00e186edcd9ae13a68a8f3030691b2ab20a8b418c6, 160'h55555555555555555555e8535cf5393398b23ce6, 160'h333333333333333333338b6537c655855b9e248a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{346, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d3cf5669d7a6aa345133a0ff9f56a88c995a340d, 168'h0094f884562ce27b0b67e0e80e486c4d4e2264e651, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h55555555555555555555e8535cf5393398b23ce6},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{347, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c2e0b6b5d370f374f3b2f5a2e4a01e2bf3c2e158, 160'h5f6879f63a40a9cacc8343214ec2925c47f1d18a, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h49249249249249249249a29098d23107a7743433},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{348, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b43dd1c55ca1a5af0e9ef4f3b3d30c70feca6f4d, 160'h4fdc2b3171e117fc3e058b7d0ba8818f977ca6d4, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h333333333333333333338b6537c655855b9e248a},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{349, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00f3be38c3aeff9324d740bc7adb0fea5eeb9ea64b, 168'h00ad0a634a2d199bd2023affd7a7546b645fd0bf78, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 168'h00ccccccccccccccccccce2d94df1956156e789229},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=168b(21B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h0a9c2a9de3f46939ef33a03a607090ef3971037d, 160'h7742033e020fc35f676fc650d170cc300deb261a, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 168'h00b6db6db6db6db6db6db816697e0d7a9322a28280},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00862e2eb41fa97389e6d9a5809f33c476255e851c, 160'h6c97ca144a98c842e706d73431d90a366dfcac6a, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h0eb020c9b97c56649802d1e8ce928dc660acbae8},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a896b2ce7de0dc53d813053a64a45053f9e6341c, 168'h008f3b7c374dc223c0ff5e32cfc517856ae25ada3e, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h55555555555555555555e8535cf5393398b23ce6},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a6b2f424d53ab1dce8ded84894b7c935daa2d869, 160'h576c5baac08c1c5ff45e2b4f5e2c743e24661c7d, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h49249249249249249249a29098d23107a7743433},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h299d0559bcd39fb4a5287989d5a02a93ea21db17, 168'h00dc64a6f176f66233d1ccb92bcdde100d39793cd4, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h333333333333333333338b6537c655855b9e248a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2d785f5990bca636e04238d50ab5e3b97c9cef0d, 160'h7d41f1eb8e50f07924c775a041567268fd4ac49f, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 168'h00ccccccccccccccccccce2d94df1956156e789229},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c0b952451eafffe6b5dee5409e8520622ae877f6, 160'h2730450893af945fe327a600458068bbe2ba2ebf, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 168'h00b6db6db6db6db6db6db816697e0d7a9322a28280},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c05720b3bd92b0f8c72bf85c0772166217234020, 168'h0083a1a12194eda0a5aa53f17f7bff65d6bf5fbb08, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h0eb020c9b97c56649802d1e8ce928dc660acbae8},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{358, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 168'h00938cf935318fdced6bc28286531733c3f03c4fee, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86, 160'h24924924924924924924d1484c691883d3ba1a19},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{359, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 168'h00938cf935318fdced6bc28286531733c3f03c4fee, 168'h00894b5a17a0c6db3c257cae09057a136f93bf9de0, 160'h24924924924924924924d1484c691883d3ba1a19},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=168b(21B), s=160b(20B)
  '{360, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h6c7306cace702312943d7d79ace8cc3b0fc35c85, 168'h0176b4a5e85f3924c3da86c3eb284543c6006dcf86, 160'h24924924924924924924d1484c691883d3ba1a19},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{361, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h6c7306cace702312943d7d79ace8cc3b0fc35c85, 168'h00894b5a17a0c6db3c257cae09057a136f93bf9de0, 160'h24924924924924924924d1484c691883d3ba1a19},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=168b(21B), s=160b(20B)
  '{362, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 168'h008c8b7f800bc9c5588b4970e7559eca926fa38e7b, 160'h6c5d8223426e1cf8d2a2791ab710a14305048ad3, 160'h2e3567b523f24421cf59dc80925775b148eb5380, 160'h38aa38f17c131f0128af4dcafe01e68305414586},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{363, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 168'h008c8b7f800bc9c5588b4970e7559eca926fa38e7b, 160'h6c5d8223426e1cf8d2a2791ab710a14305048ad3, 160'h69b9f46ded69a35ac00a053ef9dbb47d073d6729, 168'h00d059cb77081101578272ca48bf5980c5019febd5},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=168b(21B)
  '{364, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h008c8b7f800bc9c5588b4970e7559eca926fa38e7b, 160'h6c5d8223426e1cf8d2a2791ab710a14305048ad3, 168'h008e641a5d857f8c86963cace4f89537741da1a32c, 168'h009bbe6d38a198847906223f08dc6f3a8ecee563c6},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
  '{365, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 168'h008c8b7f800bc9c5588b4970e7559eca926fa38e7b, 160'h6c5d8223426e1cf8d2a2791ab710a14305048ad3, 168'h00f036a3151449a8f854c12c6fd55bd9fb02ee67af, 168'h00c3bc5227188b85b9b9c33fa7c5088f8e8e02de86}  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=168b(21B), s=168b(21B)
};
`endif // WYCHERPROOF_SECP160K1_SHA256_SV
