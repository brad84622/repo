`ifndef WYCHERPROOF_SECP224R1_SHA3256_SV
`define WYCHERPROOF_SECP224R1_SHA3256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp224r1_sha3256;

localparam int TEST_VECTORS_SECP224R1_SHA3256_NUM = 261;

ecdsa_vector_secp224r1_sha3256 test_vectors_secp224r1_sha3256 [] = '{
  '{1, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 224'h2f396442932cb80e2cca3381ebf0d975f33f6d7b77da96aefba1216a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{2, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h8ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{3, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 224'hd0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{4, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{94, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 248'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e7632640000, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=248b(31B), s=232b(29B)
  '{95, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 248'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d30000},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=248b(31B)
  '{99, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 248'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e7632640500, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=248b(31B), s=232b(29B)
  '{100, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 248'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d30500},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=248b(31B)
  '{115, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 0, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=0b(0B), s=232b(29B)
  '{116, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 0},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=0b(0B)
  '{119, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h028ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{120, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h02d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{121, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e7632e4, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{122, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb0853},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{123, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e7632, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{124, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 224'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{125, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 240'hff008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=240b(30B), s=232b(29B)
  '{126, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 240'hff00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=240b(30B)
  '{129, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{130, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{131, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h018ed6690a135a8f918c0598c2d2fee3b4ec7c59a4dd66a65b6ad25ca1, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{132, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h8ed6690a135a8f918c0598c2d300b66f2b0a7928b5ac53d0b21a0827, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{133, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hff712996f5eca5706e73fa673d2d0032edf43c9699367682e9f189cd9c, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{134, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h712996f5eca5706e73fa673d2cff4990d4f586d74a53ac2f4de5f7d9, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{135, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'hfe712996f5eca5706e73fa673d2d011c4b1383a65b229959a4952da35f, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{136, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h018ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{137, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h712996f5eca5706e73fa673d2d0032edf43c9699367682e9f189cd9c, 232'h00d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{138, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h01d0c69bbd6cd347f1d335cc7e140d53cfce327300afdfbbdbbd173310},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{139, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 224'hd0c69bbd6cd347f1d335cc7e140f268a0cc0928488256951045ede96},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{140, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'hff2f396442932cb80e2cca3381ebf1c2d312867d3d63fd6d699f44f72d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{141, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'hfe2f396442932cb80e2cca3381ebf2ac3031cd8cff5020442442e8ccf0},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{142, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 232'h01d0c69bbd6cd347f1d335cc7e140e3d2ced7982c29c02929660bb08d3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{143, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h008ed6690a135a8f918c0598c2d2ffcd120bc36966c9897d160e763264, 224'h2f396442932cb80e2cca3381ebf1c2d312867d3d63fd6d699f44f72d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{144, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{147, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{148, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{149, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{150, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{151, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{154, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{157, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{158, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{159, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{160, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{161, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{164, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{167, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{168, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{169, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{170, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{171, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=232b(29B)
  '{174, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{175, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{176, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{177, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{178, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{179, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{180, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{181, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{184, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{185, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{186, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{187, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{188, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{189, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{190, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{191, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{194, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{195, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{196, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{197, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{198, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{199, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{200, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{201, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{204, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{205, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{206, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{207, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{208, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{209, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{210, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{211, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{214, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{215, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{216, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{217, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{218, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{219, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{220, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000001},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{221, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002, 232'h00ffffffffffffffffffffffffffffffff000000000000000000000002},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{230, 1'b1, 256'hb2d2232f6d22c49f89c3c3a8a99484abbe828ffe8430eff4b891ec16ea512813, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 224'h7eb5cea4bda67eb17c42fd9e4ef8fc07a386c4d38b8e3fd7ac14e601},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{231, 1'b1, 256'h00000000713791d986ab76aa7cb5c46cf5a62351efb6c1cde74a8591d9c2fed9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ce9c8f262a8fcfbff26a2ed56156dd7fa00df1b8dd78f28522f9599f, 224'h3f8b90758650031ac943b6e89a2d401c03a4845f4825385edb0b9949},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{232, 1'b1, 256'h310000000051db6185687c0e1d43cf6f7302a7ecf3fe3d6bd30b5363dcc85614, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a596c710492f86b31d7c3031ddffa41eb6ecd0d255272777765d965c, 232'h00bc0e0d134f359088438f9d4865184a9134b22dc930a32df317cd2dad},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{233, 1'b1, 256'h80e10000000005f3acf7efe73a0182b5f719824bfa118c4925a1e8e0f194add8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h44bf0e8ef31adcf935bfdbdbffb848160ef5d5f97973303503ae43c6, 224'h58194109101107d061575d48aefb8791da1aeca9214fcc4bf9b60dec},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{234, 1'b1, 256'ha4392c0000000005c4dc1e6e2994620d6a959373e62fa5f6e84cabd790d6e56b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00bcc56b38d6a7b227a00f235f0aeef3ebf846cca2db14c29027339fc4, 224'h4355863fcc75f246f213a9b4867deb2a7face8cdf5dfbbe43f8ac31a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{235, 1'b1, 256'hd7cf0d00000000000e615ec0f55109462536b34045963901b95960c6cf5296a6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6ee3c0f02dbb1c5991fe897f8534bc9ba39e3c4a5c31d2326cebfb1c, 232'h00e85b88cc3b25e3f6c9052993d3b43fb1e0d36840c64fbfb0b979f74f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{236, 1'b1, 256'h8b9d7d14000000009051340f34c75a0e78f4a191b3f908bfdaa334f32eb47b51, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h21dd71ac10881ea88296395ab8efbe822c081b5a6d448e6e5d6de917, 224'h3b906e2910ac307a545c7c5e5a4155631be6ded9da8719f4590b5df2},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{237, 1'b1, 256'h432701b4c5000000004e77e86a34ff07f3069a9b547da784a05d7d5d950984c6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3c8dd1c1da01ca7793890cecf967aef7b3199be89973f40f132f47cc, 224'h7030a2afbf16e0200c9b5d9104009881b5667f5c991c3150d5ec0923},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{238, 1'b1, 256'hee4ea2312d5300000000f10e2378adc2459d7728a0eb1c3fa70bf25ffdfc2d9f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1bb538ffd49b566203b3390186d41052e2158bd8cabce482e2bd9cfd, 224'h2621fe8a3ebd93982e7ad1f876e354a56809f8cdaf7289c247a93509},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{239, 1'b1, 256'hb519e0108d975a00000000885c7dca69fda64d70ab959d0a99034d75dd180ce7, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0b6b5578395738451e59bc461bfc558b0ffadc75045c4298b00f9539, 216'h3147e9cdce81809e25b10531c59ae3f225c7a7681ff5135cf317bd},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=216b(27B)
  '{240, 1'b1, 256'h0ab9f26cae100d3f00000000d72de1818987a2554c6818367ae35f6d08dc2478, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00cde67578f4666789a8b77812ca4c057feee8b7cb2ac67e038292c272, 232'h00dc2dad5133d0de4d1d5f4e66c12641b0d036058382237da8c02570f8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{241, 1'b1, 256'h20069e1ea6d4dc3f640000000096664b82ba5b4b6bbef31881c2e21cb8b32bf1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fdae74f7618e26dcaea23d96aa50bf3132e2ada0ba519b0cca94e477, 232'h00d84fd4438476fd42fa02b510a88b8d66bd023c5080a54de3d3c8fc8b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{242, 1'b1, 256'h88c1ae896d5b1ee1e1280000000051e2c22d970dc99dcebfd57a35be0f5195bb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3a9c3646b7af34c502284ef0070287672dd2b59e2e60f7272d50095c, 224'h561225addbaab4b7bceba248b06dd462779bf1ee3198c2ea417ea42c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{243, 1'b1, 256'ha8dd2ff8e9ecfade5537f2000000005f36a2ec63912dc97f1b148cca8d3e986c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c4d91e546ac9dab2ccece18c49398d6342c0123149b598db9005320d, 232'h00955ada4cbd17e4975467633fffb2321f5b4acb23f4b3021a063287f8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{244, 1'b1, 256'haf52ca1d210a9ea8ae35e8fc00000000cec8a7eb3b52686105536d8fc3757f7f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2ffec2697a93f0c4c5a48bec8b15dad327b1b70017e6925fa76b683b, 224'h205dbac588cae4f0ed3b8c7b4101399ce183d38211ed22306d0cda12},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{245, 1'b1, 256'h913090d6f8bbd4e10e2ce1c5450000000016451243b9db301de24772cd781cb3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00fec15067a78ca643a53f827f56a8482c59d7e0ad38b07321d6fa9fe9, 224'h3ce7e45b31390e026b485664cbf64e39b19703c8ef7b0f2d61bfe6b6},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{246, 1'b1, 256'hc1cc5ad98460c3b9e3852479a3df00000000808b0b9e82f6ade0de221aaa7ab3, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00d57668679c06d00db112ebfd273f6aa56701b2008d77284f305201cb, 224'h21cacc0f2900debc990cf2aa52c67bb7a9d183f331a3b984d63a157d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{247, 1'b1, 256'h777e0e4f4ac2bb3050202e89f5cb690000000030c36872c4a1b6f19c1a447203, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c3c5260bed20289907b8b4fb6bd7fe69c257fe50fa84aaea7ec1ac0e, 224'h38eb78dc31766a1b038e811dbe6b80683db5c06c7d466b6f1bd44fb8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{248, 1'b1, 256'h8b15a9990c7fe432804ea9a57b1c8db8000000000033521f6cd85d48845871b4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h33efa91052f2a89dafd2b06cfa28b0c8243e3cac8246c1aea3cf4e60, 224'h41f964715dd55418a5746f91ecff15b7c6163fb94c18979cf693c21d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{249, 1'b1, 256'h2b623d836940fd3a612348a20a8d1caa00000000ad69c80f64d89f5f050714d2, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0085618ac165d6f879fd4f771c5f1a88019b04052c5f940ba052a541a5, 224'h6640f1b8db137e516f405b64aa09d31e8c1dc9ac4d5abab6f9f8760a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{250, 1'b1, 256'hbac4743859e5588409f25335619fe1c7d2000000000056aaa54240b186b1ebc1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009d1873a053a280bd698665ab4dd087be3080c2c3c3b9a2d728cc0704, 224'h734210e8416e08fdcbb3251f383928976443c559f50e7164f084c807},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{251, 1'b1, 256'h7eabb2d7d21887903ffba869f353928bd5000000002d3e45954e4b6e21fd30d0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ab1fa9ddd8f16798fd015251fd71a4add962afb6f01b00f91e42352c, 232'h009d71b11fe1a0628c012cdd938e838acbf22aebd64c1da01d5b2fbf4a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{252, 1'b1, 256'h951cd3b90eec711648999d2ca3e8e821b86c00000000574333322ca94097a491, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00869f3ec4765450ac03aa2a4a632d5f7a9603b4b52f37029dd2c7289b, 232'h00a4bd2d056fe243fd3c6d719041b2093c81125f0ee7752730c3987311},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{253, 1'b1, 256'h01ca3636d480cdce6ee63cbe3665c7bd88995f000000003f5d61628138af2b7a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0fd7a377de13b55ed9e39abed7153ab72b3864ae00089be6cb39c5ae, 224'h01999722036ba44e9e00574b3de46a7c2af46974f3ce38181cebace1},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{254, 1'b1, 256'he64458ff971279b567c8eb016ac86c39f963cbaa0000000056fbecb71ef3fd7b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h179ff07fe7b684e7231efcb22216709b6c5b64f3e2ab2b6962b7d0e2, 224'h3077af624bfa19a3df87362e3a41ea0e7f904b32c06851cee0f5b6a1},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{255, 1'b1, 256'hb15bafa66eaa8c73cedfc9568ac5a41a5b0a45e38e00000000f88ffd117bf4eb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5d6817bbbcfa633f934456ab5946744128bd0eb7c5bbe6db16e9594d, 224'h73c234f3f23187b318b984d099838ef57873ba6de48bd9fadcd2effe},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{256, 1'b1, 256'ha0daa5e1d6fb10cf91937045a9adcd668e53d8d302a8000000000223f8bb456a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00adf7cbd33018fe58d3da640dc8dcdb5db75a85b8409ef8a6d34a88df, 232'h008ae5cafe6833ad40ea2698cd862df9a5718f3b00935885f89134d9ba},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{257, 1'b1, 256'h4b28f92a09aff0587c6eb0a61588a5f2d6b1e85955436500000000ecacd385fa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ba7720511153b6b96a38635e9997caff1ac31cdea4023241d01f966c, 232'h00a0e72ea20c55bba47ee6aa7da3ebd1c1dbafee7152e3e22778644026},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{258, 1'b1, 256'h1d29293e1f2113a0eec5780d25200ee18779ad86ca0431390000000088a9c6e0, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h10a8cc92e550c816999c0a9bde2b345a2a75c6f66861f060ff2a3742, 224'h6ef54556c7883fc45e8b00638ff76c1f3eeafa895e4f2dce990249fc},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{259, 1'b1, 256'h3f466438a18ea4e57a572e3ee501d7919c87bb35179a13bc5a00000000023949, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2980c3af3b6fe6fc5f0f82e74b848453cfed1460cf99a080bd5a8566, 232'h0087d3abe0bc652743a75a54579a34b82a91c488990157c4a93645402e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{260, 1'b1, 256'haa2ef39293ec474361e7562735439b835b55d17b130df2421eb200000000fc40, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2c3d2fef2d23ea431f36dd3258127326f83aba9989754fd733931bb0, 224'h64de0f37c334eb07f57e5dcf925a7806f90f1af34c2544cf3d4d9f65},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{261, 1'b1, 256'h1df7127ff896950a28abfee5f9dd0da5da0f5960cfb1d46fc1617800000000d9, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5f08496864ba9b6b74810405fbba579a5aecca52c3c9851bce3ae580, 232'h00fad2d32d584679eb0074285f34d5ee452ed0aac2222950bc3cb01960},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{262, 1'b1, 256'h69e86af97404788bda6b6925dd727c578ada594a03d4975b545b70a800000000, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0755fbc0cb4847101118d266e826cf23fdc664bfc4b9425eeb567342, 232'h00c2fec316397cf167c1b234a7bab46c2a26b6b48b87790325995bf9a2},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{263, 1'b1, 256'hfffffffffbda4755bba6de00c2701a0c6fd32c7e4aa1d876140f979cc80f34c6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h254485afee6912f38bffae771553aaf734c779b769e792b2623ab056, 224'h6e599ea2fe87d2228992cea340b14d8872ad3cb2abf35a1f453c7c24},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{264, 1'b1, 256'h22ffffffffacfab2fac775cbddf678eac83d9fa2dcaa8379ca3af3fb8dd614df, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h0099e668983f0c3c4168081d376646074358e923b05c8be3080ed0d2a0, 232'h00e0b28c84f2ca323d89def878debd019f3a895c8deaccbe69b56c4807},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{265, 1'b1, 256'ha92dffffffff4bf463c8eca0c62afb2c35c2a592ad8e8e688aa521a258f47338, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00acda06a1f01dbcd49e8998e2727755cb6462baf32811f204351589e3, 232'h008ee9d910bb66295817c32d69b53ed6eabfa2e09fb39d46439a8a481d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{266, 1'b1, 256'hd0fab1ffffffffbf5c5a0dc94820af6ed2c80b5411be656e273b963141464e36, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5224c582ac8f7101bf6fe14a9617ca0a9878dbbe026ae230d1e63d0f, 224'h61f0e486a1b7cce228874e7ccb6dc8dc95434afe6dbb7494b9f0e1c9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{267, 1'b1, 256'hdf0ffccdffffffff58bc3fac8197329161b5dea9f0043e8cec2a9a631ea38cea, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h009d05470e3988f76e782684ffd743bbd3a2bb683b0f2cddc873ff79ed, 224'h3a1a4e796a78475db7000407279a665a2c406793110415e5655b6698},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{268, 1'b1, 256'h4d77a2c899ffffffffb8c2d8566f592706ca04276262ff7cfdba0b2ad6e2a6c4, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h74d5a5f801ab103a8de9cefe365753e5e4e24aae88b18ead08f9e7e1, 224'h22195ff2b1dff4f8ef7382a52f177a766a8f839b65b77076850c5edd},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{269, 1'b1, 256'heef9d05b88a0ffffffff18a16611a3f3ac44331426f2bdbd5af203e092e61176, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00eee00958aca3b5bc3ff48533ccdec3eb565663f173367cc95a9f314c, 232'h00ebc3ed0d610e0b9fc63d8123b927a333af6ccc2fc1404291036e514d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{270, 1'b1, 256'h7e6d3c190be6c8ffffffff27a4b129531bcb4fad150112ceeeeb8d10098dcfaa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0f0a83fbdbb05c611f6430a8d2f47c53e445831c878203cb81513878, 232'h00b4b1321f09a3ab5e4cc27befd89506651a4e40e22af69e58b3c88691},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{271, 1'b1, 256'h0edd238c04bee70affffffff0ae88780ec5271030a1847cd73f722925df9dd43, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0a67da525ab869f3c6bb4dcc1821c2ac065728cd22d49b0ba5813ba8, 232'h00b70065b12a6d2bc592783a7942ae0dae3ad1e7c6f27cacfc2b48dddb},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{272, 1'b1, 256'h4dd115320049ee2e9dffffffff0de268e472eae1699ca5afb5c838313db94bed, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b41f01a5b75fba4835798156ac882e82a2e29859960132195c1f7e91, 232'h00f421fba6d0061b92f8ab8ecbe7b5791bc43c5106c9ac9747e5da671a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{273, 1'b1, 256'h1a1109052e9ab4f5dd2cffffffffb1e4604e058f3040a4af85f1f303bd3830cb, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e3163b6dfd6585f50ac934bd25ea86065eff6376387a56cc210897de, 224'h05d93a2dee9a55228dbc3df260152c458f8dd6f72b1d57f37f6f685c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{274, 1'b1, 256'h6162159e82cf80a70b34f2ffffffff193b3c777305a8fc809337cb13014edc7a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h27a2c5db14c60f71c3f08196356ea7094db6559a4c5c7ab097aad799, 224'h755741a777ad419b5c1853bc6f8da89c282a67f71cd1fc3abfe6ef1c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{275, 1'b1, 256'hb35876d301bf4040fac24355ffffffff7fd82e02fe5885a42240d05fff5fc61b, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h6b5c4a2123721cf74e151a3f3d97880d198cd7850a490b3736ed28a4, 224'h4b0107b4c7f32a46315160b39f95d2bec469981960eeaf99f30e8d8b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{276, 1'b1, 256'hc5ae766a399aa8c082a59a4f62ffffffffab6578abad5454b86f0be4e36bedc8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h219a8f9d6701d7b51d82b293d2f0ce4847e13abe9dfe8de426164040, 224'h33623e698063becd8f28445ddb16caedfbe093a2c1d89925c28a12f9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{277, 1'b1, 256'h619548e83b2bf592724b244359f9ffffffff7ed41c49517b65795ef980c30f19, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a0676519c127f56b025695326eb68c5438b5d473c6b81b25d53793c2, 224'h62ce33315ea1ae83dc48e7e774d701dc27b364484e3133de24f08e19},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{278, 1'b1, 256'h2ca970c6acc18b4ad3b023ba01ac4bffffffff4fa0a25f4f35f9b408dd09517f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00b16cb831277a401155134fb30d6938b9918665af7e59530fcd9cc0b2, 232'h00f85a29c79b30ab6d9439eaece5901d65774ae1893ac603e3308c29ae},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{279, 1'b1, 256'hbd67ed69ca5085f9326153231b96b177ffffffffffb1a4447142406fbb23dd5c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4eb1f5dd75615bda8368b94566dfdda9d7d8917f1863d3604059fb4f, 232'h0080b5e243be6219350f60af1b50578f3d6204b5efcda10cdc338d08f7},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{280, 1'b1, 256'hacfb85a5cfe484ca5801b819b3e4159dffffffffe10cb294343a640526d5faf1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h600282c901cc3a4c8596a059b5ac217a9b999f0d3b69b24b3917d1cc, 232'h00f1f401cd8cf106992244b3674ed9e55909b8683357be44fd48a1c3eb},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{281, 1'b1, 256'h62c18f3f3271e3341a7d3033529b28a2c3ffffffff4e9cf2e8ef755e0953597f, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h54c666a30d72a0475a4cf0fe0bb58f13aadb361ffba89325c56ec48b, 232'h0091f36a9fca040343fcc29c7fed35adb9db9a2f17c1f35de4afcc8f0a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{282, 1'b1, 256'h2df78ec6d8628aeba725a007584b63636883ffffffff0ca2480cb4e3523b2daa, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ffea346481a37d7f2728e2bbe35083bcbace7b91e06da2ad1825dbdf, 224'h06cf6eee77ea7a4da0ed79a8a167adec51c8a2de906f3f7fecde799e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{283, 1'b1, 256'h07fc58409c7cb5c7169a63d09e4de5120132b8ffffffff1f95f5e389535720ac, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h38fa40a57e4a04024c899051cc8080c5261dde66ea59fe532e852013, 224'h3e99d123e596e993d677683bd25889549155edae098e59a29fe7d9cf},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{284, 1'b1, 256'h383dfba6e0aa10f820e15e27374c2eb6996baf43ffffffff66a94ff532236f85, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7f62a985c5bbde0e11e0250a97d73fa38011bb83b6fa2d9836bf5c45, 224'h3bd850832cc305e6b7d9566d36951ac4794b2d08ff712b18b0af6594},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{285, 1'b1, 256'hc41a8affa1bbbe99587538b31e0b61f8b56ebe58d7ffffffff45e1ee3efb6c66, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h311f063576c8373b96cc1652ab3be3a58eadea786e75b17a04c2bca0, 232'h00bdb7096d675d1024291702dd991d5606c125e6129554922e02444fb1},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{286, 1'b1, 256'h26fa9d690a2129917bc3520b913f913f1f081bea9aa3ffffffff0fd642c24a4a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h65db63a663e35fb97ea8f0752a3190134102f4fbbedd14bb5c1349a8, 232'h00abdfe68c7f0c674f302488bc030558d35649f9a9c69d5801a575cb0b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{287, 1'b1, 256'hb291bf1a8c66adc9def9a0a96da478aa1d09e06797adcdffffffff8fb0460842, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h075ceeeaa2ffbe5dc173d84df71145a056500a90f8fb902a24c0d363, 224'h688cefcf26f584f8d598da2b960a512b6b65a425ed536a4bd570cf83},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{288, 1'b1, 256'h81d64896fa11ee94e49755c0180cc0478de87bf9969ae759ffffffffb4b7f4f5, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00f84074b42b14acb8715ab229e4261c09b096a58b69f510f5f491ba6e, 224'h304fe4129c6dbe481cc92d9dcbea983e40eafef17ea46039608a1431},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{289, 1'b1, 256'h3b88244a6ae111bc752afc8f997cc9ed1f9d4079a0f644f3d8ffffffffa41c42, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00ada080ecff37ca818f48dd5c0ebab78a645e973e138435637237f870, 224'h4d85eb195089c83c92b483a53b036b33050aa14ba244eb48a0f97d9d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{290, 1'b1, 256'hbae669421b6378571d97fee160d401bf8f4698bcfa6788a85be7ffffffff6844, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00a7c22c1d68e8bd563520cfc749d7de43d9ae045187a2424168eaacf3, 224'h6959ae2c1fe30b45b049c4a5e418654711f21cbb925dce89e51a9ae4},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{291, 1'b1, 256'h1f52ed3bbbeeaa23026b261a17bc00058f2e37cba29772831b7ed9ffffffff02, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2ce15f3bc4f827e2cd5f59b7980f694e91c4b6a7b77c616f17121136, 224'h3f71766ac9e52b98f58a6895112e43b75925183a29a73bd835f95593},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{292, 1'b1, 256'habacfdf5c9518bfcd685890b4e11728fe6bb738a9517baacd701149affffffff, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00e69b6b3c9a08da2a90d59ac5454c10246bd8dec06590420391140693, 224'h52d090e54b79fa780b46000a070b1a78ba9797b34b1761f09408c80b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{293, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 232'h00c1a527a3efe3b397bef889b699b192a7663d9d60449dd9eccbfa8e55, 224'h7ba2de0347d0895c6a24b26e80044586f6718beeabc316f18c88f014},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{294, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h008e761a8fb0ae0f4d077c8331039186bacafac74ad25c499787d09ef4, 232'h00af5e802921def07b85dbaca11146382cc4121767d8cd0f0798e2bc0a, 120'h00e95c1f470fc1ec22d6baa3a3d5c1, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=120b(15B), s=232b(29B)
  '{295, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h008e761a8fb0ae0f4d077c8331039186bacafac74ad25c499787d09ef4, 232'h00af5e802921def07b85dbaca11146382cc4121767d8cd0f0798e2bc0a, 232'h00fffffffffffffffffffffffffffffffefffffffffffffffffffffffe, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{296, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ca50630a872adcd558c388ca3b024cb59e1299bd45d9e324f605e261, 224'h3c69a70c60f49e04b38e3738c5e591edaa51d7974de9e72725d8a690, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3c, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a3b},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{297, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h1977aac0b91c2b65f580a5f33d8045a3a56e3a3ab48d8613f3ac0844, 232'h00c315f37b48cb771635e16afbca84948b9e4e35690a0990bddc6cab9a, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{298, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h041ed3f4d372c3b7c4274e15c1a4c2e52011a5ea686de23b3b27bf3f, 224'h6d8d6ebfa63b7467a691d6da259d932ece80b6ba946d992ca78c3aab, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 232'h00bf19ab4d3ebf5a1a49d765909308daa88c2b7be3969db552ea30562b},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{299, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h6731bd2f7969febf93fa2382bd4fdc93ddeede8f2deac4c3abf1ce7a, 224'h19516b15727d111c786b39ba11026d25a220b4fe52c5f56fd4ca5dec, 8'h03, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4aa4667eacd6788f17ebde59e78dde177b2b378945ba487d325567d8, 224'h5d887d32e8cf6d5182433d8f81c945b4356d3ebc0e970dd0a9035387, 8'h03, 8'h03},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h0322435ef8557da9306c645a0b614c6f6ce98d859697784cf74f2f23, 232'h00a8cd9e243e9088170133bd81eb6cd28571fcf207509819f443e5bbb5, 8'h03, 8'h04},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{302, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h0322435ef8557da9306c645a0b614c6f6ce98d859697784cf74f2f23, 232'h00a8cd9e243e9088170133bd81eb6cd28571fcf207509819f443e5bbb5, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c2a40, 8'h04},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=8b(1B)
  '{303, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h5719bd78776367ffea95b9313ec825c70a3252326aa1ec66bc207bd3, 224'h327ae05556f62f5650db898b316e689b5c377a8a64d743a89ab4153b, 8'h03, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c6f00c4},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=232b(29B)
  '{304, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00bb1e97c4b5bedec0af97169db06d040647bd40fa7853c8e8d0ad430b, 224'h1025ec677e900574853cc5ce761a92bae929ec86076acc4859beacc8, 16'h0100, 232'h00c993264c993264c993264c99326411d2e55b3214a8d67528812a55ab},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{305, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b00ff7e1925b9717903a05d40ce9860ed12ebed8c686e05a9205a976, 224'h110ee94a9a3267ab1565c66cdd5ed2844ccc5c6a7e78e4821b954f98, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{306, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b4f18d031097f179effad146f5fa7e8574e6493dc4133a7e6bff6763, 232'h00b11ad9abcde8a93b78b6bc1f71d96168712263f6fdeb1da9b1193912, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{307, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00a35240c68e8f4ecec640ad2cc54533275cd6b54f480476e0412f191e, 224'h7c4bdef2aa2561fbb2d26f9034836265b81e555d56b6f446b6b863a8, 16'h0100, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=16b(2B), s=232b(29B)
  '{308, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ef67cfa95eba7f21e47e9f80e624d06297e3c516b5d4810bc03264f4, 224'h7ae076453ed06bc43999b713aafd0eb2aa8192f61a61d6560d66a3d8, 104'h062522bbd3ecbe7c39e93e7c24, 232'h00d05434abacd859ed74185e75b751c6d9f60c7921dacfbb8e19cdba8e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=104b(13B), s=232b(29B)
  '{309, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ff16dbdd1335d3d31acd1fea3cbdd5fafbcfb13367cc5831574a0bae, 232'h0081763ffbd6bc8720d46e7ee3cda01b98a0cf479816ea46bea8aae199, 232'h00ffffffffffffffffffffffffffff16a2e0b8f03e13dd29455c5c29bd, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{310, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h009c88d34bcdc70a09bd9cb4aab4e40fa900472d635c4ebd2366e5d4b9, 232'h00ecc54c3d44714953766bbb1257a3580a2aa85170e418969ba3a66841, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{311, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h009c88d34bcdc70a09bd9cb4aab4e40fa900472d635c4ebd2366e5d4b9, 232'h00ecc54c3d44714953766bbb1257a3580a2aa85170e418969ba3a66841, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{312, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00a3ce180bd65ffc76d5502ae806a6b434d7e69b39b1940e44c83604cb, 224'h4150ca512dddf3363897dd8d23f76564412188cc9be77c170dcef4e7, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{313, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h7a1183e83dd8e38b2aef19c9e604a205ecf50abc9ad1b2bf3a062ba9, 224'h35d0ec70d1c66ba124872a47d044b8bb7b6a405b9a9bcce636f9e788, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{314, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h6fbbbfa60d49b603fbc7f6f6c922df0364c03f089af3a288ce4337d5, 224'h28c46eb6f43e9c4f2664ff72d587cd706c620cd718bceb1197482ed9, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{315, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00d50a93a475ab04521ca4bc4dcd06872e85fc587a7c56e68a6e94846a, 224'h4511f0bd21af19dff4def09b04bcb20e21ad21e0f8c4a49f21856aa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf7},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{316, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4a0298d7a7a670d2538f6aae65ddf6be35d474bbdd1b6aa0a812d974, 232'h009251866f630eda71e9d727964e563a2596ec04c4d0134fb997021ca3, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00a8ce483b42fb3461047c96ca00d0c226ee2850b79192346c7ce37d46},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{317, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4a8ead5e32234b2a78171bbe3215f1b721f9ae113c7e9711bd44cb28, 224'h15580cc1e9f22a432e8070f700b949ea55cfcd9323589fe1edb06053, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{318, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h55bd003333e449dc59e181cb2e14e2240f26bc7f3f1713a73ba0e36c, 224'h69ac8b1fb9c4c270ec57a6afd3f8c65f1e34c5176c7f7684e861167d, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 232'h00aaaaaaaaaaaaaaaaaaaaaaaaaaaa0f17407b4ad40d3e1b8392e81c29},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{319, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h7036b96d9033ea5bf6a63bc308936da1636b22c601f5fd1a3fc8b491, 224'h028417ad37899b3ea1dca7b67ec60a7e7b0af04d024bad8aa3a5e4a3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00c7bb3d419456ee8a53d67867550ed5eb3c00d55638ac6d2132bb007b},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{320, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h58fe2f40f6b361167bd9757e73908b21a8f43c420e13aef119211e64, 224'h6775a49681e2d646dea26bf257f8f7fac9f7fb2e9bbfd36649957b84, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00aab6daa4628852ca4b25e917ef4771547c75d5ec5127c9c6678cde4d},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{321, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ae5524a4533101a5cfe3907d706cafa7f904d9dfe38ceec59457d62e, 224'h18434e271edf58008c15d627dabbf5691e9c9eaa7930094ce885e2ce, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h008063db16787011a1c1212af044599a91f78869bd790f5dc588d842e5},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{322, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00e0af4ad4f06a41c72d502d6934c8c3f4b34f062d1cf723b3712c9af3, 224'h4a3d09ffd3506e11669609ea8fe8ee54b30188bc0ad136cdcf73038c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h17688246313d0b42a8ce483b42fb1f0a6217394611f2b177ada94b47},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{323, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00deaf785750eef0b3e178ec726956b9338838b0be79ca5166041937b5, 232'h00a6b69318efc4961a50b44cd4b792c271539f3b4129e8e8dadc9684b3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0088246313d0b42a8ce483b42fb345942d2565666e25fd2f85a60ebae2},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{324, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00e14fb7fc849de20d33c6c5e6b358f5ba702eb2b9121def8d3deddbdf, 224'h58153c8e0ef0b78993f4d17405c1fe2b20880d40b229f7de51a4d6b3, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h1048c627a1685519c907685f668c11b76a11dc9e381d35c5efc14b87},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{325, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00f83a254c07c29022454c43be9bd5e99c630ff7d83206713a1fbfa0fa, 224'h017a0adb068fb28a9418328eac1bc19c6c92c3f1666a773250571a19, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h313d0b42a8ce483b42fb3461047c69e7886089d9f0c0fc2c4d917952},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h23ac1ccb807f76fa99207af67f662fb1ee10f1d5fddb715eafa8ad3d, 232'h00b18eceeb7432c70250f8e92fa990baab18296547fb7901acdd8faf59, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h1c22615f35d488bad614c3cc5578205bd25c0d73ed985e1214d094e1},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{327, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h119d9f0c5f5f6206df598622ec7afc756a0c1c1b3d1133528a7a06cd, 224'h0df17a9164719714488b9ba8021885d4eaa83e8842b11af368d06304, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3844c2be6ba91175ac298798aaf040b7a4b81ae7db30bc2429a129c2},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{328, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h008888ae9b1ab8d57b18468a2c16f8c971a70711c6361a9afe14be4e33, 232'h00af32311a18ef6b965c8f6e252051794a3467de9f58c06a8545b743dc, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h5467241da17d9a30823e4b65006861137714285bc8c91a363e71bea3},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{329, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h2ce5a3f2b3fc7916953ebe71a7ff33921cb57167abaa871a07202196, 232'h00ea2d3b61820bdd5264f060680844d7217a21601e3ed37a79d5953b98, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00c031ed8b3c3808d0e0909578222c589a6c20acfdc6764385729a3691},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{330, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00bae5f11eb77e354a0d0e33c4ce24839d726e1700e514ccbdede23145, 224'h4ffd009fbeea9c7307938f8adfed84de3600920286281d267c88609a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{331, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00d153ad8f462d2f9388fa8b43517aa2a7799dea0bbb1fba67c5674172, 232'h00df03b778b587abc18db23bd52f43913714d1f41b8c91907b24cf1ef8, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00855f5b2dc8e46ec428a593f73219cf65dae793e8346e30cc3701309c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{332, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h39b30cf6827e95c4bb1cf5a201e3611ea87660c671fcfe4837a55ba8, 232'h00bf990d7e7756ab4c0f08f0d674980caa2e559c93c84f7042fbf0ace0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{333, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ce72f433416794d9ba0e53735eb2277ffdfe84f852ff06b26b2ba48d, 232'h00cef033d6f897ce820f3178f0331b475ad9f8e6be2ff34788e09e55c4, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0084a6c7513e5f48c07fffffffffff8713f3cba1293e4f3e95597fe6bd},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{334, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h69211fb68e0ce40b590bdfb262753d3817a9777cbcc18292f63d9446, 224'h7fc0dcf4d6a02a0daf952f1bdc99ecb4bcefde8d7eb22ae14be44b5f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{335, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eae4a3d43da31e5bbb6767ec18b03c22314dcde77f6adae7e6a1b66c, 224'h3b2b6f2abe22f00376703cda54a6b6e4cbd7bac7614782ef9e94b26f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00d8ea27cbe9180fffffffffffffff3a43fa3662a899627950d4eb64bc},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{336, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h1a51969a30f966894ed0e1b763da7cdd2a258a9a9d6efb019419c152, 232'h00fd8982295489e97f2d8d6ebe0409d759a5ca25cf9627f20e39f1e651, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{337, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00909bb6c47b981b1eb3ad78d6ad6b04791f9952429f98a01416b778fd, 224'h6c38107d55d28e37493d22e2aa2a4c66c9da2cc90be2202278870f92, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h00bfffffffffffffffffffffffffff3d87bb44c833bb384d0f224ccdde},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{338, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00eec9dbb6fe5ed5c8e4f8309cd81d506005efd52dca73e8874957db2c, 232'h00840f6693e77f92088c6e411075ff15817ca0f6e669a295d01d2442bd, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{339, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00a4b5e9304fb04bc6257fed45083fc7f50aacffb962d42b3b3a6c6177, 224'h58aa38fe0aa034025e4b7ed045eea3edad0a5ece26bfa7441239f521, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h7fef8ed425081537adbe4773037d77ccec1a3dae490c46360c92d067, 232'h00e5309792680df204f3ccaf51d9e73543f21e519377b504885b6e55c5, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 232'h0096dafb0d7540b93b5790327082635cd8895e1e799d5d19f92b594056},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{341, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00d4c38c0df6f7743e577ce3d054a32e84b2a7418d1a9e00a0a1d30e13, 224'h5428f7047f7eee01b2377ac2eb041d24637f40977b11b24f2904d9dc, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h21cdafc19b3c56e71933d3692d76c92c00cd08d146b2ed4c03525393},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{342, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00d4c38c0df6f7743e577ce3d054a32e84b2a7418d1a9e00a0a1d30e13, 232'h00abd708fb808111fe4dc8853d14fbe2da9c80bf6884ee4db0d6fb2625, 232'h00c44503dae85dd5210780f02928b3d927171c578f8603d16b240663c7, 224'h21cdafc19b3c56e71933d3692d76c92c00cd08d146b2ed4c03525393},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{343, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ebc69137db89c0189696ee75ff03706b0d939639bb64e220d70ecee6, 224'h23a446d65b083da18cb14cb6a9e57f007558386065726ea34feab573, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{344, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ff8f64c0c0f7f0e81d205b67a1c3bccf0c3dcf3bfdfdc80a61471e80, 232'h00a0cbbf29ebedf5381016937ad91335c5801bbe6fd4a1ee6199295601, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{345, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h11c0f94fc2820ead7b14208d0620a35f376f1c10b6af16060454b048, 232'h00b004d5322db3039c7fdd4888fdc0caffae81edbe53e80cd05df210b9, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{346, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h3e4fa16464ba762f06e7cec2fcbf66269ff742c10a53361217f2053e, 224'h706b308fa36b5de586523d32244eea63a4d86f215930eae2bf99808e, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{347, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4825b311ea6b6ad86eb6f8fe9d29eead7a7a93daafaffae356a785b4, 224'h73160b436b4894f5ee3f50288dbdb66fe1c08f94f677ecdc5eee6e44, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{348, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h235c610afcdc0a22f84d753b1f7b9cee388f8f5d68127046500b4f1a, 224'h605e49168429c44e190d3612f355bd7e63978fb6c9a61dcd53b13821, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{349, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h009f77906d353c1b862ec4794687c69fa506405c4d0b57f4ef8491dba7, 232'h00ce9e810af65edf1ae583e6f9d6f2ddbc01365e1e744f2987af5527e0, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{350, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h31699a0079058d604ed7f87c9aeb44bf1978527bfe01025a0cdd2a0b, 232'h00eb919883753f880b47d06a1acccdf7d77bf984fa48f26c959b12fe7a, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{351, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h3ffe7230477fe2ba4c3fd54ab1da6fe0c29eaa5b6c18982eb7038a2f, 224'h3911699ad8e6c713a7ddb2c7d569f1ae648b1400115e416b2be74c36, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00db6db6db6db6db6db6db6db6db6ceed4c09e84c77ebd9116e17391eb},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{352, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4abf00bb45592cbfde38b5381d1847bd8816d9113a99b18b7d1a0e07, 224'h1f47d0c50e5506c06af9e4db68ad58818fff05df0116048a0418b951, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{353, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h17564764dde6c5d5bc1ff0cc65478522aa0492cca7ecde374e5019ec, 232'h00c17e0cd326b5a30a5131097da640ea1f81b577ea98df9e5906574361, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00cccccccccccccccccccccccccccc121be6fa59cb431754377d168831},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{354, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00ad728313f562dc2284a6f6c4a102c569c3bc730279248b15d75df168, 224'h0e900506b8e46beb36600bf2e2a0bdda494dfe3fbb4221b4587938d6, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{355, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h38b185b1b7d7497db0ebb1f0998575706bdcc0c6b4301c5c99083210, 232'h00ea4d43854b92d8c3aba8163803893095f448fd6beccf5ba90e6d075e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{356, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{357, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 232'h00a8ce483b42fb3461047c96ca00d0c226ee2850b79192346c7ce37d46, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{358, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf7, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{359, 1'b0, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 232'h00a8ce483b42fb3461047c96ca00d0c226ee2850b79192346c7ce37d46, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{360, 1'b1, 256'ha7ffc6f8bf1ed76651c14756a061d662f580ff4de43b49fa82d80a4b80f8434a, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h2a8e4fc8c813be0459fe6fd5a449fcd27118121180f37f96857498fb, 224'h487fabaabee79f667da6505c5c171d299732d37784fd73775dfd3db3},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{361, 1'b1, 256'h5a7a8ec92299354caa012069a923d56d0043b22408fb36ff8cd0ecba3aacb0a4, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h1e5a15190a1d2631f2222d704489041f72e0c50548fd526eda975e1f, 232'h00ebff8dcb8c1134ac5dfb271182495590fc8fd8ea7b0a4f7f8ec78900},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{362, 1'b1, 256'h5731b7c4bd04cb9efb836935ff2e547bf2909f86824af4d8df78acf76d7b3d4e, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h295e399cbf4904e22850240598e009d6b40d6391e370aba5a04042d9, 224'h2a0c5841560271a38c7b7c3bb064990e204bae693e2171a246942d40},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{363, 1'b1, 256'hf3683c9e3da9a7f90397767215345efe3be07565f14ab80d102f50644b98fbfa, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 232'h00f04e2dc4d8f01de69a5bae38d0869be1926e0ca75a641f2fcd7784d7, 232'h009613012233db115ba180f7363aafbde09dc0a5ebb6707613838a1413},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{364, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h4007008e430202f9577e43a0b21ffd169c046d5bf35c2b530115a618, 232'h00d845d27c3ab6d1f81881f1c5f980d1c25844a484a87c99058d76e3b5},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{365, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 232'h00917e785e5e0432f597d10dc400725a0344cf4856be31390573a1eaf3, 232'h00b85d30901195e05cbef0e282a079f5c229eae8eb282be9176df9ed88},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{366, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h3e4f9883f7acaadf2a076234fa99fd25a5d8369fb7766aa5b2eb3fd2, 224'h42cb3e2eb9f5431fca4a7ec83637aca92fbebe8afa4ab4bced1088b9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{367, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00f33a24a2cd64f41d981ffa97c24cb73d28379146824c8d4c77c37f68, 224'h7019a27bc87ab06d3a312b3027215104044ab9a917de5542071a5702},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{368, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00ff961228b94551c201bb61c15286d119e02db2f45cdc66979debb3a1, 224'h34a490221e2bf3097d369f3fcf9c6507a56780051f54ff961f773e20},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{369, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 232'h00ddced52bca9640b1a1a7f85bb12d8cf36f0cd60b27ecddd2a944dc49, 232'h00826b3c1a839da54a8beeece69da8681c643fec79394d982dbf0c6837},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=232b(29B)
  '{370, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00d8f0e29a424ba0a53ddcb8f48fc4b65019d01e7e8dac3ff63847dcd3, 224'h62ec0f1f7b36512ee98cae1fac6bae7505e84e6eb279623e064fa094},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{371, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 232'h00f5df25249adba5717354fea143b93793f32ea8ba31cd377f9bbb6eea, 224'h61376f02d5e7517f1cd2a5c36c452a76decb282daebfeea5a5b32e12},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{372, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h4b9b6fefe18c73272ee66ab96fe340b3835b1f63f903b1ac76ba3457, 224'h0c580a65c53b48d1180f0985fe0f9d5f57cf7eb5e572b9714411aa98},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{373, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h6f72f5934d17a126d0d6fe0afa599588c51963023ce93c312ec77baf, 232'h00d5b4b96943f585cd1568a617e7c47b9dfaddfb58bec13c57c15a0a10},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{374, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h1579cbc71f2c067d1449c5eaf32e121eca057a35f375bdc93f771a3c, 232'h00c5e865acd21b480a65150e7010e5072cc5aac16e3316fa8fd32a078f},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=232b(29B)
  '{375, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 232'h00ee501caf390634fc3757ead8e3f62e5c8e86c0448289ae5dffc6a30f, 224'h36d39f3560c5afa05787248787235e8edd8c42e713ed43adfb82879a},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=232b(29B), s=224b(28B)
  '{376, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h714796f7fe64f4de33bdd8eaeff4e7e3a8ea9664a0d3249e07bdec4f, 232'h00ec82e64e1c6f652d1198c2996f893222d920d36d7e38507e86f37357},  // lens: hash=256b(32B), x=224b(28B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{377, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00b010d489c9661c1a283537428868c4b5bb29d9503de697ac574d22fd, 232'h00ec677ca1c8b12eb0304cf090d952c63801ed9c82d751dbd76d4bc18a},  // lens: hash=256b(32B), x=224b(28B), y=192b(24B), r=232b(29B), s=232b(29B)
  '{378, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 232'h00a8fb6a1a558cb2221560204babedf6c44d48109ebae78d27e784056b, 224'h1e532d50e0b6721e9345248fcc37593077c4bab575b55d216fa2a3f2},  // lens: hash=256b(32B), x=224b(28B), y=192b(24B), r=232b(29B), s=224b(28B)
  '{379, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 232'h008085d6b7f3d979356f2a213bb243746ea678e96a705e6893bf2a51f7, 232'h00b4d8be5c3f996ed40af1024b3a8c9f65c90efb41d8c5987aca115524},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{380, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h5f1adbfcde7a0a929f43ba30e0d88ea2ada5b4a8bbf55336eb228fdf, 232'h00eac90d6f0679bdeefc4284027c5e527cab4cb27619217783fb2c421e},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{381, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h17b20a24457e94f8b882a4fc99692c2c44b5c853b9c234d03ad473b3, 232'h00b03bf47ea4533e86229b96c65265423f89daadb9f3f69b0ee37c21bf},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{382, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h00faccc9c38ebfa8e2748d32f8c41cc291c4a2b27cad4a411e5119d19b, 224'h70e5ba90a65e03515594c919f17eac4d809596e6a2735b617b3852ab},  // lens: hash=256b(32B), x=200b(25B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{383, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 232'h008f8e90c2a830534593bdf1e5614ed9ca75f8253956d17579a6a4532d, 232'h00800c2d43eea0b7211f739f4e75ca5677ea0efb109b094aac354af676},  // lens: hash=256b(32B), x=200b(25B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{384, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h2728cc303c3ed54a05a371f16add7c2da6d2277b80a932b7b9749df7, 232'h00ad2c93f83723c19e20385fab9116188114a1280be7d1fd9a661e5e77},  // lens: hash=256b(32B), x=200b(25B), y=232b(29B), r=224b(28B), s=232b(29B)
  '{385, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h3a224d4baaa5d5c332a3d62043b1aaf66b029880010c839c5c033aa3, 224'h2de87b37b0305cf6112e0ac94200118ff493c0a379f4beb0b6602e02},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{386, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h009159aa74a88b5917809605e14736a00e92f4aacda2b87dde950a5ff8, 224'h4bd456c6914cf21c88be0bc9c64a3d0d7b2cbd5c776297fea3a12f5e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{387, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 232'h008b21ed26d9455613a0431edb41d4227fc5711d1a6c70e4e0de801737, 224'h2592becb967e25d234a2516986c18a1c687b2969db7178cd204d30c0},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=224b(28B)
  '{388, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h5c7c63a63a69787bfc469ab70a6856f7f322447f9ce74573d0f94d2d, 224'h3e80ff0a9fbd8c11a08d7dc02237e435838de2d2b51eec1156e667d1},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{389, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h036b3f33ccc347d6f0ae2b9e79ef85351d06e61870b1cb08054c909d, 232'h009a27fe9d699cf6e2c2ed2ed70c9692f1f6b96fc5b4e50d9926a752ad},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{390, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h3131bcf930d1136df1436c4780c095e00170cecb929f6ee71c7458f7, 232'h00a1c6f0f97cad156078d248fc7e7974045d27888e8f6528af66047faf},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=224b(28B), s=232b(29B)
  '{391, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h1023fa4d5dcedab53a8fdfe2a8f8da941be08c63146e4ba2ed87bd4d, 224'h367a88e393fd1ee4ec925f7f920d4c3fe3ba48edbd253261ec706c5e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{392, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h00b525fb6204d3d60fd406b1066f0ae4bd7ec75b0adfd807de8201f10a, 232'h00faed757f5a68d8a8338788ea531d6f7c85a88c9a8bae7f696ebb6eba},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
  '{393, 1'b1, 256'hf567a849061ea8289d35c676e297544ec6d13169498da7ec0ed827f1899ce6b5, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 232'h00e472e504ef4b293b7f4a6cc99ba33a702f35593f49cb284137776b44, 232'h00c1efe440463fde3b604d48319e0ddb93261ae608d009942a01933241}  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=232b(29B), s=232b(29B)
};
`endif
