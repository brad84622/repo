`ifndef WYCHERPROOF_SECP192R1_SHA256_SV
`define WYCHERPROOF_SECP192R1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;
  logic [511:0]  hash;
  logic [527:0]  x;
  logic [527:0]  y;
  logic [527:0]  r;
  logic [527:0]  s;
} ecdsa_vector_secp192r1_sha256;

localparam int TEST_VECTORS_SECP192R1_SHA256_NUM = 231;

ecdsa_vector_secp192r1_sha256 test_vectors_secp192r1_sha256 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'h508423e042b52945e2198ae8b4a97d3810961d886c6ce1e4},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'haf7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{3, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{96, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 208'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a030000, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=208b(26B), s=200b(25B)
  '{97, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 216'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d0000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=216b(27B)
  '{101, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 208'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a030500, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=208b(26B), s=200b(25B)
  '{102, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 216'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d0500},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=216b(27B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 0, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=0b(0B), s=200b(25B)
  '{118, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 0},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=0b(0B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h1a4abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h02af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a83, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac29486546cd},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 184'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=184b(23B), s=200b(25B)
  '{126, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 184'h4abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=184b(23B), s=200b(25B)
  '{127, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac29486546},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{128, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 32968'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a030000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=32968b(4121B), s=200b(25B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'hff184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 208'hff00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=208b(26B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=8b(1B)
  '{135, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 32976'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=32976b(4122B)
  '{136, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h01184abdfc6df2ed2d0c9c706749344af637f86e5c3461b234, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'hff184abdfc6df2ed2d0c9c706815765a8a0f20daf8cabd61d2, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{138, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'he7b54203920d12d2f3638f9850aaad3fdc735b55807075fd, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00e7b54203920d12d2f3638f97ea89a575f0df250735429e2e, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{140, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'hfee7b54203920d12d2f3638f98b6cbb509c80791a3cb9e4dcc, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{141, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h01184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{142, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00e7b54203920d12d2f3638f9850aaad3fdc735b55807075fd, 200'h00af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{143, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h01af7bdc1fbd4ad6ba1de675167f147334184175dafd376e7e},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'haf7bdc1fbd4ad6ba1de675174b5682c7ef69e27793931e1c},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'hff508423e042b52945e2198ae91aca8501fc2a53d6b79ab9b3},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'hfe508423e042b52945e2198ae980eb8ccbe7be8a2502c89182},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 200'h01af7bdc1fbd4ad6ba1de67516e5357afe03d5ac294865464d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{148, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h184abdfc6df2ed2d0c9c7067af5552c0238ca4aa7f8f8a03, 192'h508423e042b52945e2198ae91aca8501fc2a53d6b79ab9b3},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{149, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{153, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h00, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{159, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{163, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'h01, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{169, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{174, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{175, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{176, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 8'hff, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{179, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{180, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{181, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{182, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{183, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{184, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{189, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{190, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{191, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{192, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{193, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{194, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{195, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{196, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{199, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{200, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{201, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{202, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{203, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{204, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{205, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{206, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{209, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{210, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{211, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{212, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{213, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{214, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{215, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{216, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{219, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{220, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{221, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 8'hff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{222, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22831},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{223, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{224, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22832},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{225, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 200'h00fffffffffffffffffffffffffffffffeffffffffffffffff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{226, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ffffffffffffffffffffffffffffffff0000000000000000, 200'h00ffffffffffffffffffffffffffffffff0000000000000000},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{238, 1'b1, 256'hec8293d735c00c63847a99e43f08c510d279009ec01e5350b0d56cb8f19465ea, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ca3c599e99ded921130f3a1afd34dad6b0f02efd13a8df17, 192'h12c9cb2405eb711785a3add143b054f3cd74499a2bf916d3},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{239, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h6f20676c0d04fc40ea55d5702f798355787363a91e97a7e5, 200'h009d1c8c171b2b02e7d791c204c17cea4cf556a2034288885b},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{240, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h5c6683cf0b0867ba1f80a3c83a740c6b25d067a15524210a, 200'h00c9ec84d890fd8457598d06be72984f6384291b2bd98a9fcc},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{241, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h1c1af41c461fd2e7ac90cf03775430863e0625609392d689, 192'h56621316c3fb0fc17d1e140c87a8d25141ead133b66fb543},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{242, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00837f82d3e38cc20ea4e8fd37cf22b3fe186f5db7887fc9dd, 200'h00c91f2bad58385cc572cf4c5eeb6ecd57c07c55ae54eadbf8},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{243, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00c9059b71d8fa9fd88a098fcc8af33b9f80285a7bcffda023, 200'h00c8b24dd67c8bbb00d05ba9a5d5d7883b1fc26dd1cb6bc385},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{244, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h1eba3835f014e1c0173cd60a053fadc9fc0e7709919496a1, 192'h64c7d823cd73423b2c7966c0b248a65e53aaf80af0ab2b50},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{245, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00c788e831bd1cfb700034e72f65d0bae19f9466626515e302, 192'h7c9bf5755f2c036c3f5f771796c41c7852f30ac4e1d58307},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{246, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00b50ee502ffa2bb07dd0051094918e80daba2021acfeaa536, 192'h48fc394f05a742002ac474ab27d718babb931fd031bb1afb},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{247, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00c0e6a3260f71c47914a52fa2a982805837a266fd57df5a48, 192'h5c7cb80e4c7724de8c35b754b49ff98af83dc6a2f9fabd00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{248, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h0081a675a2534f28433bdf9c934406b70d38d95fbf292afac2, 200'h00965a681f046b676e7983ccf795ac1d48373a76e5309de6f8},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{249, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h54a5508f5d8244d34ccc5fe0d964ed2cce612aa602ba8bb9, 200'h00fb9e8253241677989c6cf51edf16b1d48375520df7043ea2},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{250, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h230b4df715ebfe839ced490130c89037757c89a2715c19ef, 200'h0088c8726f7a303f507ba2d767ac727b6b673cee1588c87818},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{251, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h008c8dba2b4c277168c65aa9398e63f2098e4bd52b07f57ba3, 192'h629818c1e0c4c99a23148b2c42fe568ef0a5e2b05bc375ea},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{252, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00c58940187da3be8462df9db7bcb3d8dbe0415f6edc1b5f93, 192'h4d92f7377656b962327564e2261221b270c58249ef12ae54},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{253, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00cd59fab71c72b0cf8e22a3b311715505c55bc9ec0b629a34, 200'h0096d877ba0cdecb45eef4bdad96074ce09349d6f6fa09d049},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{254, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h125b39558823f19874183fc6193c50e4f5fd7f87561f43b3, 192'h1b164d656157ee6fd5c6ed20276f2f9e8e78f40056f4c917},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{255, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h0d7edccdad3379dcc50513397b2988ce4f200f08363a21fb, 200'h009bce1635c8a59bb79b6e75b6f90ce154d4375bf8ea54c2ed},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{256, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h008d043f335315f492005b55d0b9ce7b622d4a57ce546d41ba, 192'h718ebcadc80a765adfae660c2dc14627da4046e5b0757493},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{257, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00f9c31b588329bf386d30eec4e18eda4a6fa80331cdab7fd3, 200'h00839015b1c469d077791138027a18f9cf95c1f6c26038fd9f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{258, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h4d23bfb770d8b60bb7ab1aa45e1f6b1da414945fd52215bb, 192'h2d2c57ee3fc517793470f61f38e1ac5dc9cd88618d7f2782},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{259, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h3f5ec831bcc1862a106a455c6342ca0e5a16dd87716f34a3, 200'h009f586b8cd559ee0aa4c2aee2ea7085e86fa94aa2cd439b98},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{260, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h424d505066afc412387b147f0cf96e1ebae3a16f0c0d69ef, 192'h446975a09f8d9c20d2704196f1446f354e79ff3d308c7e48},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{261, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00ff310f50a988062a42c214906af6bbe8f16401e6d5f2feb2, 200'h00b6d48aea808b89082ef8236554b7d08001ca9e9e75f3a46e},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{262, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00c92fa70af822dbc54446db3a14991f1b1a259431404e74f9, 192'h3943d5a2a8466551ec71c134c8ab3898beeee8ebcc515e57},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{263, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00d39ba286b249286df48695023150b201f340e8e9b2f8d841, 200'h00d1ddbcda01e59a13b82e601d8f0c377e6e16c23e64d6c7d0},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{264, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h31cdf0bf4b77c10f5f11bb2ab2a3c778059e076824146523, 192'h058c3be3e7d01be17f1d135745d581ccfcf03ae0ab6226f9},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{265, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00cb5e28b4704e678dbc176d29e69d6ac0faac007dc5bd1eff, 200'h00f5aeb3cb95f35804e14df45e6560d15883c703cd6b6d323e},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{266, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h0088cd865f89d4c5188b8e31340648ecca5090029815f317a5, 192'h5442c7016eb2cdafc25d90923ef3c8a2d7c5a8bc56b6dc61},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{267, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h0a666bbd50d32922eceb07fd63971d6b44c06e39f6ae37ce, 192'h13df79819941a6413a4f3ef6f1b62882ecc88b30b041e3ea},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{268, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h654c558777a4fa29fc22026156220258986a262ac65dd8ee, 192'h608e8dc90e569b3d182a663e93f740ebc9fc7b9cd5112879},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{269, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h3247b2b9f8f59df93efea88267609d8a8f7c45a216a2ee20, 192'h4212ee42824f30fafce4fe8286b69cbac02192fcee13e32d},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{270, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h37479876e1e96c7ad149ec7725e07ec16ce30f4a849d2471, 192'h1dc2e3642b717b8d1b73b9cf94d8ff070c0b7eed4141f0ff},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{271, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00dc12856e8545a1b99e3078c41311a76a4d2153b277b2a5f6, 200'h00a5562129d77b60ee20cdd96380d169eb227e47d62ce8a792},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{272, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00fc441581f33e606b1eca2243e677369fb9ac94825d999af4, 192'h72d505027448b937a5fadfff6fa21778459d7a090e68410b},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{273, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h5968579514668883386e05d6d5813f8e3ad54ab595fb51a6, 192'h35006e924c80a145666bb097b9ccf6bfa1650d7b005869e8},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{274, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h0086d113f6cbfcba4f4d58dd9e0166ff6f6c317f24d57d53b9, 192'h6c0a580d47544cb58feae35dac2437171b02a4eecb306801},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{275, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00a644bedf78ffae253536f3e6d2cceac8878f7fc037b8316a, 200'h00b6869fcce992f506109ddd9ac9124e911b27d56f2bb30e27},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{276, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h193f5680cb656c321307f0cf016c3647d9daba2fdf847f79, 192'h167304e7d677d139103edbf6d09a4291aecb6e05719158b9},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{277, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h008fbfd696c501e6f7feaa971e80691466907cfefcc1a96ef0, 200'h00c6fa2a35bc8cebdc4dfd70262bf0c0a8bb4addb4f3c17bc8},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{278, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h008b3bcaba24580ecaa8e730a29008f825a2f683bc3b314d10, 192'h480e092be161b4874b605b69a23d6b971b7205c1da76c56f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{279, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00819c51c1c3e9d65b7eb26718f50d3673a1783492af6c6403, 200'h00b3ebd329221b9022c4548b1b73f590be3659d8f89fcb63d4},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{280, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00db0a95bb7c3fcd6193d712a6fb9002c8649b397faea4a3a2, 192'h3a0144aa631bb232eb937502b8f5e7c351d449d6807ad50b},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{281, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h15cf54f4362efcbdce3a559aff7e2e1307614a7aeba25b4d, 200'h00fcf2bea5d38678e60b0d0df55116212fb9b4bb1013c5b4f5},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{282, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h009d4069399d4d8aad19b31f33cbbaff6a614cdde3b11496a9, 200'h00bed1eec79772b64b8014f72a66f5152ba0de5eaec72249a4},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{283, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h4f720842ca4677b1c3f54f5800f328b37b420fdad97b4c82, 200'h00befb5c561acacd99c88e851f07499765ff80b9384b971ca2},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{284, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h0bcc3e54ac1b14c1962d86204a9bea9fb8d2e4b3b6cd7472, 200'h00cfe0b094b669c155e32edc03de153482d5bda6428712d243},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{285, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00e6c02360d53c1b870af823685432a0c9d92f7ef4f5831c82, 192'h230399616677856165f7ec24d98a7d1a71fb546c735ebc65},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{286, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00a30170d6c1518c766d91b8be2fa1c9527adb075417480204, 192'h4011aa3fb5b3ed22f5567fa52103bf992df4962c10d0872c},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{287, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h008cc4670ec57cd542d4d355a12949d072cfb0dc38426c62c6, 192'h033e389e84e76211db83dae6fb772dddf50ebf544832e042},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{288, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h634dbc50a74338fe4d0e187111eb776f88a2b7034b879dab, 192'h4201e22c4a85b3232f21ed346ac335e069b610163fdff242},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{289, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h33596110e8d4a1b6c49d3d619dc24c153bee63aed3c35778, 200'h00b991c1bfd346ea8013696aa29711a6bb7ceaa5050d074521},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{290, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00f560fe32f05e37c39c1b96c1ce6629ec8d9774acba0a2dec, 200'h00d4c008e3299158c83bd925d540a8137697f791532d5be5d7},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{291, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h314da19b75e5f8116ab7c6a671e7dadb379a8e86c7452c7d, 192'h6cd48d19c8667db383385742ede00007e484825f214065aa},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{292, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 200'h00f1bbe301dd0a1e766b58bf812fb53808bac91e6f84ad9e21, 192'h687352d26ff14b2fc1fd5f18ffccf9020898b6fe0419dba2},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{293, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00cd35a0b18eeb8fcd87ff019780012828745f046e785deba2, 200'h008150de1be6cb4376523006beff30ff09b4049125ced29723, 192'h6bec819bb205c55575ddb4b30022a04886d6d562e38ffc22, 200'h00a9cf7350956fa86fc9fc7703388453df3b24bc0e4c5f0be3},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{294, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00b02ebfa6d8365f7bf0d1f19a0fa407eb4feaaa7dfff8675b, 192'h341b88c93b0be1173fade7befc78aefd0847e862b13f32dc, 96'h662107c8eb94364e4b2dd7cd, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d2282e},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=96b(12B), s=200b(25B)
  '{295, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00b02ebfa6d8365f7bf0d1f19a0fa407eb4feaaa7dfff8675b, 192'h341b88c93b0be1173fade7befc78aefd0847e862b13f32dc, 200'h00fffffffffffffffffffffffffffffffefffffffffffffffe, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d2282e},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{296, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h1c2bb4254256a329ec973fff79951c895a53441f2b73e4e2, 192'h5daf0bd36c2e64e44d0e517b49464cec34daef9699829d22, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22830, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d2282f},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c422742cb5d7f990dc9579e85a0339da7ecabda11d7d18eb, 200'h00f547da5ec37681ce86916fc7ef4e91b76aa2073f17531cc9, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h73e5f9eaf96c8c84c93bd31bf65daf4ed20ea0ef67ae0bd2},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e70f06da0e6036bb0ee47fe47836a0f4382e3349ff927112, 192'h6feeb50ab0f618a5557e488bace8fa2932fb03009ed622a0, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h41a92de5298636d693e86db59b3ed26215e70ecfe43620d9},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0094e936a4149ababae26300ec4c915409f6bbcbbce94611d3, 192'h5f326034990f7993559d97901e7ed1808587378cdb236c07, 8'h02, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00bb41507556b67368feb9978e7879305e4fa81beb2c95ad95, 192'h5d7f0e5c3966ad5fee2b5901cc3dec4190175246935ca993, 8'h02, 8'h02},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7e18073ab95a26038e5f35a805c76c8b880f9d175793005e, 200'h008be399eddfdce76e1a42ba16d065bc7186c08b32fcafdfea, 8'h02, 8'h03},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=8b(1B), s=8b(1B)
  '{302, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7e18073ab95a26038e5f35a805c76c8b880f9d175793005e, 200'h008be399eddfdce76e1a42ba16d065bc7186c08b32fcafdfea, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d22833, 8'h03},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h29dfd732d3c13161364d2987d312c9308b8a1dc8b4f05dd2, 200'h00e5b139e112b780fb34ba03903a6c23e7691627c6d6f07e82, 8'h02, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4e4feb8},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=8b(1B), s=200b(25B)
  '{304, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009017d4ad62933e72336feacc1bead950a83089de8250a794, 192'h00812bb07b9991cb9b5143feda006523f8570cf01df138f4, 16'h0100, 200'h00c58b162c58b162c58b162c586293ddc4f185918f2cca7bbd},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=16b(2B), s=200b(25B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0095e29b80d6943da6e053dc1e6bb29180a3260d0e055aedd3, 192'h2ef8f9f432d773c0ac7ce51f51868ecd4ed3745d9baba447, 56'h2d9b4d347952cd, 200'h009776c260bd6a78d36f5e21dbeb71c84d9d1dd348d5c29843},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=56b(7B), s=200b(25B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009e89eef90b6c71347513445c3edd12b921f5eaa249851213, 192'h6be9f9603e3126de833ed6f760d07d5a87eadb2095135028, 104'h1033e67e37b32b445580bf4efc, 200'h00bd42bd42bd42bd42bd42bd4271c1ba7da5827d34af84755f},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=104b(13B), s=200b(25B)
  '{307, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e8e4a8087fbb956cb784d2cfbbd4fb10fc5b82dc52992132, 200'h00bfcfdb9d6a4079b70212a9a547f165673441cfea068b86f7, 16'h0100, 200'h009ea14637a98e63d3c3368641e12310b8fae991b42b894a70},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=16b(2B), s=200b(25B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00a5e0079778dfcc1546f4f3b7071032db86681e32aa110698, 192'h094c333ea7f796eddc157607828019414f0641b321c3d288, 104'h062522bbd3ecbe7c39e93e7c24, 200'h009ea14637a98e63d3c3368641e12310b8fae991b42b894a70},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=104b(13B), s=200b(25B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h138e1036185e32e26f24ed6e747c92bc5750d3b1181d20bf, 192'h1abc97cc3f9f648bcf4ed10b6c8a74100bc9c18460de7e5a, 200'h00ffffffffffffffffffffffff99def836146bc9b1b4d227b1, 200'h00aaaaaaaaaaaaaaaaaaaaaaaa6694a57962f28676788c1acb},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=200b(25B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ebb8328e0c8bac41eaf502dfb9e5f5d57014c7ea842b6617, 200'h00c7b6fb10434359da7a29ae458bf2b03b7c9290f79c4196fc, 192'h555555555555555555555555334a52bcb179433b3c460d68, 8'h01},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=8b(1B)
  '{311, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ebb8328e0c8bac41eaf502dfb9e5f5d57014c7ea842b6617, 200'h00c7b6fb10434359da7a29ae458bf2b03b7c9290f79c4196fc, 192'h555555555555555555555555334a52bcb179433b3c460d68, 8'h00},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=8b(1B)
  '{312, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h73761b8c8aa66d47c302a1af56ce6e64c139de565a2de1ec, 200'h00a526726d7552e162df2c42a7e1523083e150be83167c334f, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691418, 192'h555555555555555555555555334a52bcb179433b3c460d65},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{313, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d7bc9b50e8bff4bb2c6c8116a25a973e95717fd857fad573, 192'h3eb089b00237660aa485016da2f6c3bdec88cc1cdb28eb56, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691419, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691418},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d02ae497238e2def130607b98eed7693a2f8ad4f9294e3cd, 192'h5d8fed9551ff73ffe0d3877cd364ffb104690052cbd0f7e2, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691419, 192'h7fffffffffffffffffffffffccef7c1b0a35e4d8da691419},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{315, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d5e7ec9b4724ad94507666e9b1e4763ad17372537966090f, 200'h00840633cdab3497984e5f5d36eb8e2a0c048a73a10e0893ea, 192'h555555555555555555555555334a52bcb179433b3c460d64, 200'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c88},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4f9a2b948e4ea950a2ec9dfda5ad1b9b619f9eb678b27cd1, 200'h00aff08eaa1b956963e6af3d61f2c5812ce50145fdfe74c2a3, 192'h555555555555555555555555334a52bcb179433b3c460d64, 192'h44a5ad0bd0636d9e12bc9e0a05bc56531434e1ee89ab1ba9},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4dc27b674729ea276d1f9c9b031f2db841497db7ce50845f, 192'h71838b5b21bfb0b238ea9e209ff89c88f8d070933d7f5531, 192'h555555555555555555555555334a52bcb179433b3c460d64, 192'h555555555555555555555555334a52bcb179433b3c460d64},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c3b346d4066a2528aed586a999462aed82cfb361aef75a08, 192'h7578d73662260bc96ca5c09b8ee279f9701a196a45c002d4, 192'h555555555555555555555555334a52bcb179433b3c460d64, 200'h00aaaaaaaaaaaaaaaaaaaaaaaa6694a57962f28676788c1acd},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00af7cee273d57a8393cb468e561a25f8ba08699cecf0ac932, 200'h00a6490421d495caad3773466249d5e547922bcf18322ce89c, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00e91e1ba6ba898620a46bcb5197f5861a6304d3b786ee744e},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00f05d260d24704880c60febfda3e2873e3e45a412d264aae5, 192'h5a4c5eaaeea3a2c8f03b2feba6a3d5b0a84f9b8538de9f39, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h0094cedff8715e3845c128caece9832c826ac733817b6560d5},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5a6289c4fb18c344a4edcfd89105c62ffa20cba6814e74b9, 200'h00fd11db2d30eb3b9edaaaead049e57868be475208052a0da6, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h68e686f0eccb840bb80bf08e2ee70d64264fd5162fe2159c},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00d916e677f68e917c53565a6761ca655e6a31ed2270314207, 200'h0094596ff9667203d4f167aa5c022d758b2ee2db538591d0c5, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00b587d583e05abb0744a5ad0b87f7e2831bce821bd28e21b9},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e8955850e22d5c08c319b66b9abf74387fe6d209356b671e, 192'h3cf26e4a6a6df3ccf2aeb15a3d949d382a7ef87cbbc419ca, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h7d583e05abb0744a5ad0bd0604d88c454169c54db223a428},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h3bc30c3d86767b9896a1b0cf644b375c548a6501adc5d837, 192'h4a27f48e68f8c6546b9d0285fbaa03a72c0e0e32ec55bd51, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00fab07c0b5760e894b5a17a0c09b1188a82d38a9b64474850},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00f883e2274d25974c468bfd5d42ab28811fae32c39ab69acd, 200'h008a492829cc6e3851f9bd433a2e27d9362af718ec5c1c2d22, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00e05abb0744a5ad0bd0636d9db93b84ffaf061f18c62da9ed},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00ac3b619c03c378e6018281e70138fb656d9e79c14287c223, 200'h00d7368c53015b87e03dd88499556ab89406e5928f90094395, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h4f1696d5ba25729655f53877ae5a3c4631776eb4bad5d13f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{327, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5f4d9383af8b02db95e63e4ac6f2e89d0736af3a8e5b2358, 192'h434b4b5682b944d11707c012945beecf85b583a15e554e53, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h0084e74337b374d0f901569d92cd585db34282d069e43e7180},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4aa98d13e19db5763a37085a905db0c12bf649fd4ed80972, 192'h021cd9adcd2ad111b5a71f20ec343f1ae610a6ad9d9d13fb, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h008b70f22ca2bb3cefadca1a56cde43528e2e95fd5f15aee0a},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00caf74fab27fbaf4c4a1da037583d7c3ac651df9863d4c4fb, 192'h21d54ffcdb5c2cc0790c712de4d889febcdb49fe890315d3, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h16e1e459457679df5b9434ae01e9721bb166f5fa2de3b3e3},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00e1e2889b4bfed1c564391f9b1596f17e07277547087c5571, 192'h3f093730dee0a334cd63df6d31abdd0ee709805ca0da5731, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00a252d685e831b6cf095e4f04cfcda744945055d01f3ea1ed},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h3f0635d2d1dc63d37a911bb0b5c4afea9fe2a6f8243ab27d, 192'h6178cda8f95d86e2f8927ce903ebad88e944a07ed8ab3417, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h347343787665c205dc05f847177386b21327ea8b17f10ace},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{332, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00bb9315dcd7175cad8205fe853524f2c1dc5a94437d5c248e, 200'h00809d06e4fd4d94055a2a0e380c097060a19ea8aa7c0c6afc, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00d55555555555555555555555113f50240d9d31212336c575},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h6db7e7cfd64693b3826e1e055af1d64add5228ad394030df, 192'h275aa157c486b6f0460a36ec009c2c395f81dbfe3bcbabc1, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00fd4f8adcc9f7c93ada2ad4f881a7308d23c58e079dfccb5a},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{334, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c106249e39105763784d762b8daabb8443035db71c208a93, 200'h00a8b212435b6a4f18efc1036dc31a344fc48a5ab9bd4a8098, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00a3a94e7536336832484b60537103f19846b5e18f86a28b1f},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{335, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h03b643a6e4f8f8ef055824811c9625e4e7fcc13cc376de30, 200'h00dd4b194796868bdca47d7c7c096a83761578de4006519447, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h009873561529936d8c7fffffffc32e60321281988de09afa45},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c36e6fa900dacbbcb6aaca3aa6efc49b453b1bd4b04ce158, 192'h2e351f235b2f2f66a9383597c10fb311572f011f52bc0902, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h3561529936d8c7ffffffffffeab455eb8a9a41f7f1676529},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{337, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h2de010ef4508cd806b145061f5be2986c12fd98431f403ea, 192'h71037bc5d2d3d3e686518cfc719bd2c00b19027e7f3880f5, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h6ac2a5326db18fffffffffffd568abd7153483efe2ceca52},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0080ed329fcdf36f7f8a33ca2bb65a71f52864d75435b0e7cf, 192'h790c28f5a4e82c9ed3a3845799ee4dc6426cca1322db7d3c, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h29936d8c7fffffffffffffffef69e514dfd0b9ad6b3f3dfb},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{339, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h3b32883de0323161da30414ad7c5e0a771e33d71bf8f0289, 192'h67990bce37618bb3938ee9cb9c142cfc85cb148b7f72668d, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00d11111111111111111111110bbf58a93776ae3cfd26add3a},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{340, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00f30d6a74f4148d42f8f3ed364a5783032206f6bb702bf170, 192'h35f9670800e4b64a2d35ca16b6739d80f7ca1d17c2569a94, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00bfffffffffffffffffffffffafc179e159301e79573768b9},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009e74033763a653ee1eb69584268de7012905f003869a52ae, 200'h00f47afc4fb2fa6a3f1572f165ffe998e40ed5125b83f51a5c, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h155555555555555555555555444fd40903674c4848cdb15e},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{342, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h31d49b617bbd70c6177bbdf7bd7d48c4b04d3033ee2428c8, 200'h00f9032538ef821c03f6cb6891742eebfad72d45fce55fd5e8, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h2aaaaaaaaaaaaaaaaaaaaaaa889fa81206ce9890919b62bc},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{343, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c1f93e227ce3ee8dd56a70e8825b2494c244e1c7c5876e10, 192'h185684cbaf96e3a47302319971ddb1cf52073dc0a2324565, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 192'h3fffffffffffffffffffffffccef7c1b0a35e4d8da69141a},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{344, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c68987d692739b2866d4182375d205e6d2e8b2cbd438b4fa, 192'h6df95d919b1421ef9d2d74a337211f9f17b9516438432eb0, 192'h7ffffffffffffffffffffffffffffffffffffffffffffffd, 200'h00d1d4a73a9b19b4192425b029857174e72d90d5a09dba59a8},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{345, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0245ee12b35d21d485df220ada6b91180d9246c8be5ad048, 192'h58062250a1d3aaea5924432e390a5de4ffc63fc9e9641269, 200'h008738d6eee2154b64f449eceefe526444f3918d3a01281e39, 192'h4758ab667e2ea3df3455aefc647da7cc50369cef0881724c},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{346, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h0245ee12b35d21d485df220ada6b91180d9246c8be5ad048, 200'h00a7f9ddaf5e2c5515a6dbbcd1c6f5a21a0039c036169bed96, 200'h008738d6eee2154b64f449eceefe526444f3918d3a01281e39, 192'h4758ab667e2ea3df3455aefc647da7cc50369cef0881724c},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{347, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0098764a1282d3a1efd6e412e205a226a52c91200ff6728f76, 192'h712f8b75ef23d945288be4b6af16d1e22fd42bb8a8ff64a6, 8'h01, 192'h555555555555555555555555334a52bcb179433b3c460d65},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=8b(1B), s=192b(24B)
  '{348, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00b785873f9994c332b86084c86bc22ba3685a6e61fd449887, 200'h00f99a7e2167eba442af9e1080d29a9bf3b1db9a37facbaa7b, 200'h01000000000000000000000000000000000000000000000000, 192'h3333333333333333333333331ec631a46a7bf5238a906e70},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{349, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h009826be07a2fb115616e96e29a35f663c45aa6aa44acc0d2d, 200'h00ba68408829c30e55b035719117565d40e3ea8ddd656faa01, 192'h555555555555555555555555334a52bcb179433b3c460d65, 192'h3333333333333333333333331ec631a46a7bf5238a906e70},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{350, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h0093505b76fc287e7e7f0471dd11bd711305434328369d5da8, 192'h707e666839f4436ee449da037844690bbc08654383427ae1, 200'h00dafebf5828783f2ad35534631588a3f629a70fb16982a888, 192'h555555555555555555555555334a52bcb179433b3c460d65},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h5bedc2bf4bd50787b08ed6bcd1725203e66d06113b86978c, 200'h00bd6839e704b81c29deaee3a43f84e585ba4267245590785d, 200'h00dafebf5828783f2ad35534631588a3f629a70fb16982a888, 200'h0092492492492492492492492457ed201ee719058a1e2ef265},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4e95cf828614dd5192832fd2b2dcd3a734a02a25101bc34a, 192'h2055117adc6de5203c44f6dde9273320a6b76d6dd69fb8bc, 200'h00dafebf5828783f2ad35534631588a3f629a70fb16982a888, 192'h3333333333333333333333331ec631a46a7bf5238a906e70},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00c3c80a17d7817c9977c793085f3079a475eebf6197c214fa, 200'h0090881282fc0004b15eac50cebcfb189a2dcd8019865af563, 200'h00dafebf5828783f2ad35534631588a3f629a70fb16982a888, 200'h00cccccccccccccccccccccccc7b18c691a9efd48e2a41b9c1},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=200b(25B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h4023272107d16deefa43666bddecc8ac713b66ca241c27ff, 200'h00af953cafe341df8e1132f790fe3dceccb46ccca9f1da8af0, 200'h00dafebf5828783f2ad35534631588a3f629a70fb16982a888, 192'h6db6db6db6db6db6db6db6db41f1d8172d52c42796a335cc},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00f6e1b3cc1e90235e443de82a4ba54d3d530525efab707602, 200'h0084764307c6c40d056dfe5322521203770e6e73bf544203c9, 200'h00dafebf5828783f2ad35534631588a3f629a70fb16982a888, 192'h0eb10e5af0643b62b86dc5451543e9035e00a5276c1f7a3e},  // lens: hash=256b(32B), x=200b(25B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00eced81c0c456fc3238d08f92238962778b85bb596b27768a, 192'h14b06921bb4656b7e800d4cf98d06f5b381b8aa0d7fa7ad4, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h555555555555555555555555334a52bcb179433b3c460d65},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h037fe0b5d37b77b283dc320af66f7b6a5636211ccf3db7c5, 192'h09bbee2333ba7c3c8983f1dbf1ccd6dc8616459c6190ba38, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 200'h0092492492492492492492492457ed201ee719058a1e2ef265},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h37697388bfe2dafa44b03111fd3f9de97664e109edd25f76, 192'h59445a4f6e038cf3f541250ca40a89ce7d3692c9fc0e0975, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h3333333333333333333333331ec631a46a7bf5238a906e70},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h714dabf7b0ebb34a591454255c8d3435f850c35972b51c95, 192'h28ce0e186e12fa73a58572f3098914211cac4a222da1faab, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 200'h00cccccccccccccccccccccccc7b18c691a9efd48e2a41b9c1},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=200b(25B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 200'h00dfa930300cdc9ee289effdcc06c26f332b6a0ef598428495, 192'h4c2e5626703904f5643dc693062c71995e789f9c9663e8b6, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h6db6db6db6db6db6db6db6db41f1d8172d52c42796a335cc},  // lens: hash=256b(32B), x=200b(25B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{361, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h7bff39306ffc5cc10f34609435ec21eab7a3b49967f7f3b3, 192'h6c0b9346b2c981d59f77079c8f53923c496c73f7ad7d07b1, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h0eb10e5af0643b62b86dc5451543e9035e00a5276c1f7a3e},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{362, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h07192b95ffc8da78631011ed6b24cdd573f977a11e794811, 200'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c88, 192'h24924924924924924924924915fb4807b9c64162878bbc99},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=200b(25B), s=192b(24B)
  '{363, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 192'h07192b95ffc8da78631011ed6b24cdd573f977a11e794811, 192'h44a5ad0bd0636d9e12bc9e0a05bc56531434e1ee89ab1ba9, 192'h24924924924924924924924915fb4807b9c64162878bbc99},  // lens: hash=256b(32B), x=192b(24B), y=192b(24B), r=192b(24B), s=192b(24B)
  '{364, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 200'h00f8e6d46a003725879cefee1294db32298c06885ee186b7ee, 200'h00bb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c88, 192'h24924924924924924924924915fb4807b9c64162878bbc99},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{365, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h188da80eb03090f67cbf20eb43a18800f4ff0afd82ff1012, 200'h00f8e6d46a003725879cefee1294db32298c06885ee186b7ee, 192'h44a5ad0bd0636d9e12bc9e0a05bc56531434e1ee89ab1ba9, 192'h24924924924924924924924915fb4807b9c64162878bbc99},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{366, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 192'h2a551b5a39771e436de636d6259ba6afb1afa5d4d897ccf8, 200'h00bca9a6ea5d92d656c4ba4f2dd85c9d86d0e2445fd5db8692, 200'h00e71a129d6448d62998efe3978fc988213eca13b5566717a4, 192'h3d126426794e418914e5670c75a197fbd93b91d55c16abde},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
  '{367, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 192'h2a551b5a39771e436de636d6259ba6afb1afa5d4d897ccf8, 200'h00bca9a6ea5d92d656c4ba4f2dd85c9d86d0e2445fd5db8692, 192'h1c5298437de413483c777e1133e62d5b81848747b89480bb, 192'h03b56152e323216bd9d9e403c8cd229a68014f6e2b69015d},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=192b(24B)
  '{368, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 192'h2a551b5a39771e436de636d6259ba6afb1afa5d4d897ccf8, 200'h00bca9a6ea5d92d656c4ba4f2dd85c9d86d0e2445fd5db8692, 192'h497b0b598aa3559d6d415fd46c6c3f20fcfb838017e2fc33, 200'h00c8ba739cd63ac91b4dd518b6b52020ef3df72b5c366ea9fd},  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=192b(24B), s=200b(25B)
  '{369, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 192'h2a551b5a39771e436de636d6259ba6afb1afa5d4d897ccf8, 200'h00bca9a6ea5d92d656c4ba4f2dd85c9d86d0e2445fd5db8692, 200'h0091cd55bb1984e9d793f9a17bd516aa7aa597569d29622250, 192'h3996aa1d58df66bddd4aaf70964775198137c819c9e6b88e}  // lens: hash=256b(32B), x=192b(24B), y=200b(25B), r=200b(25B), s=192b(24B)
};
`endif
