`ifndef WYCHERPROOF_SECP224K1_SHA256_V1_SV
`define WYCHERPROOF_SECP224K1_SHA256_V1_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224k1_sha256_v1;

localparam int TEST_VECTORS_SECP224K1_SHA256_V1_NUM = 68;

ecdsa_vector_secp224k1_sha256_v1 test_vectors_secp224k1_sha256_v1 [] = '{
  '{5, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 224'h3fc04f62221710b2a8510cc9cdc437a622fc0dca8509d7bde7e55ce5},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{6, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 224'hc03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba5512},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{147, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 224'h00c03fb09ddde8ef4d57aef336323da542aff053ba45e6d1b38eba55},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h241b54acec345f866a6bc2c44014c0cfa5cb2bb9c8f70557c7db0078, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{169, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h00, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{177, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{178, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{179, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'h01, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{185, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{187, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 8'hff, 8'hff},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h7c0828d863ce6d6913b1c286f73953e4ae012e848a052e82afda0530, 224'h0d7e7befa3c03caaad5d76afa887f1e90a46458074f3655268994f0a},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{302, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h5e0d4c378d083719d87502c5d37d173169143d3caefa1fbe9e0c0de2, 224'h6e64b7656ac29958a7ca2b83ae97504ac97b4fe7f79cbed87ee43f51},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{308, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h6d53edf91ce58bdd92e12e2d8f55d7637edd7ee59ac6e78381ebeec3, 224'h6d5a0743de3e5cad36e8894aa07a5a07a714370051b692361ad3debc},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{314, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h6a9c1de2cb1969901f38ab2e521a5a4c2d054db43851f2a175f6712e, 224'h40d588366e72441ebf1b1cb2e3516dd500b3322f7ec9771c3d0eb849},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{316, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h5d4dbf8017a04f12d9502e63718677d241cf46cfca25413c38f38f62, 224'h077cd018618cfa428887d8cf9cc49085a7ef963b8fd01d5aaaf862a6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{317, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h1a2c2331eb8f97daf2157042ac472119bc45d661fec664483a1fc81e, 224'h305c423b008045a4f5dc1bbdd0bb7b29dcd29cd389e52a4a7ed5ac27},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{322, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h593d30711700976c78bb617a2029d0b433af7b8f706856ca1248ba27, 224'h07ea97204b37184d723520069e83c27e53142a67bc9e68e777c50072},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{323, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h49285c90a8738e3092fbf78819f5b562c7da020e4881e01fd0b6824e, 224'h33044f586ac7ecdb506e1ce3f3a1abafbb44951565367c8070541369},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{327, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h3408da6225d974875437816e5c9aa7f2dcae06b42da3d03ff92f94ce, 224'h5201beea5fdbcbfff8082937c32d95ed1a9b89121c2ed94097d73f07},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{328, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h4b375c050402389b8c7e60ff896b3ec60951b7714a7a0f89d754558f, 224'h6b1a9669881f83d75229d3cfbc4efd8d86c2d3ab2e2e8bcbcfae844c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{330, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h2bf7cc09a7405cc9ff20028aa246322acb9d05ed979c5f67dc0522ca, 224'h64cfb2076f0773e5a0a89d81a2bac2dccf2341e0f82f8d6dd23ea425},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{339, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h5cfdcd39f1a1cb8c259323823896c23f25d3354fdbad446d51006673, 224'h0bef5f32aa56df10f062d33b5e8408a9c1281c002c8f325242a62861},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h06b9c9328ee02d7828eb73697dd41de06619cb0581f16d6d224d0491, 224'h0431999d333bd4ee2bff37ce9094cf33e72696456122e11bff431482},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{348, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 224'h28aa93c8c9c2d81b7e5a466f01be0a0aa3ebee2197abff4d11edb00c, 224'h6b7d6594c1def5d4701e9875f25b80176e7ef5cbc51da250a702d65c, 224'h45373e696c28f8d2e869e51c5ba9a8e76dc04015f479e49fa354b626, 224'h6a1f35a36ec1a1d032b48dc98f711d247459d9148d61a9a6a6884d0a},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h0626c8135926a2ebca46bdba2a88c99ddab5367f06ffe11ff9c58dac, 224'h296491e4e37f21f84e28993dd0e0896cf56fa05ed411ce670d74257c, 120'h01dce8d2ec6184caf0a972769fcc86, 120'h01dce8d2ec6184caf0a972769fcc85},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=120b(15B), s=120b(15B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e65c9ff5718ade2472f6a60a0932455772d6c6dc17a0fdb9dae48bca, 224'h29d6f9569efae6aedb8380a8bc8075b04eb4491edde3514af5bd129d, 40'h0100001a92, 224'h6b40cfab3ff22bd6ef6f2b1a28398acd590fadc0b1c3d530f69e2736},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{355, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00968402f95fd321c0cf75f78edbd2f8c836f2d8b55952b820f7a0ba34, 224'h354db2bda50b742a03d972b9063f455ab0f6cf6dab448b33f540f922, 40'h0100001a92, 224'h40e62110de4b8ede6ab17d2f8ac1bce1b3230f4bb3c676b2caa9150c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{356, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2f874521547c06dbcb5dd575632a45cbac3ccc69e59ccef1a1652afa, 232'h00f014b8c953ffd4e3f157130293b0cab1739a9542543a36e90b35177a, 8'h02, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c48a1d6cc5f68b379f875e4971723299b28089019afd67628e3a6bf7, 224'h09c63f963d2656bf864e080cda07cc5d30e8f4ac61bb6ea2d5646b0b, 8'h02, 8'h02},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{358, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00db7a161f1cf83a215b43ab283deea50bf2dabf29d38277ae826f14b4, 232'h00f6c231b0fbc035998fd72431475d0c1c7ecae43aa2366f3afdf5d50b, 8'h02, 8'h03},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{359, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b621d2678163deaa6fa425ec3f7a3936ce24bc71737bad547668c500, 232'h008a6d3abcd5c6ebdf88fb90b0ff3da086b41f2df5f33df5b50b9ae879, 8'h04, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{360, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d263f43fca0fda72b3f6bb521e1bba6d50f392b81b6eeb7312a21fbc, 232'h00e95f160949fa569352497e88c56f7232f204f1aade752d8b3f21663d, 8'h04, 8'h03},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{361, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0092064e58faac9017d5fd40dacfa4da86459156c8876780a993dc8351, 232'h00ce6a6c3786b87deba14855118156f0a9af09fe82999e81f2dd46e0b6, 8'h04, 8'h04},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{362, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008a5913b8da46091e1f3521703a129057582c16c60b781353f0c2b3c1, 224'h028c5efb2add74557d0f17df2795ee6f374482473a3b7b0904f6b147, 8'h04, 8'h05},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{366, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0092f0088eff3b24fd6cfb8d99adcbfebb873c3b15fad012214d22d64c, 224'h0b7b8a94a75b60f7bb4130ccc01297c7a250091d78df6a04c3cda624, 56'h2d9b4d347952cc, 224'h0135fa9cb663a24b634b6c650b61ea744182b35e059463d8479f4057},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{367, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c9d1d50e5a5efc6d387beb9fc7aa8a73fd7597e7f2b49c8174556239, 224'h37f6d59c22426d5d6be3c0ce305f80bb8f912faf9dfe9ad843128ba1, 104'h1033e67e37b32b445580bf4efb, 224'h19e619e619e619e619e619e619e64a257fec15d1aaf17fb5d03bfc17},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=104b(13B), s=224b(28B)
  '{370, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00fc64cb84f8f635864a29fec2897e8be844e54839d8f20c028b0f4ed1, 232'h00d1a9f5ebb38cfd8a9449a90a6dfbd73faf9c60a440919ab56e5dcd10, 120'h01dce8d2ec6184caf0a972769fcc0b, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b52},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=120b(15B), s=224b(28B)
  '{371, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00ca0b442aad1e1d57c43c67d7a648797f344233537b8dae6ddd248d5d, 232'h00e3994babccac8782cc18e56ce18772a2add8ec4d47fb807756390877, 72'h009c44febf31c3594d, 72'h00839ed28247c2b06b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=72b(9B), s=72b(9B)
  '{372, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00f39dc37388cb4c34fe5d5a1f2aa6041c4c108ccc13e42c61f0c418de, 232'h00adb51ba0d123842cbf2a83a8a75e2a3d2bed11adf11784d15278c550, 104'h09df8b682430beef6f5fd7c7cd, 104'h0fd0a62e13778f4222a0d61c8a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=104b(13B)
  '{373, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c8b6ea8c530305db5ad07d53d51d61858a13d2bf766541040e7acecf, 232'h00f255573d8521b52299bdcbf2ca5cdd4e00bb14dec6a07b7df5a56e41, 136'h008a598e563a89f526c32ebec8de26367a, 136'h0084f633e2042630e99dd0f1e16f7a04bf},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=136b(17B), s=136b(17B)
  '{374, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h49f6f1d2a600142eaaf7410097c1a644a91349fe8677963892d68c86, 232'h00a0dbf7abeb84ac9b5b2129b4b7e4baad0989c990321f33e5edf1ced2, 168'h00aa6eeb5823f7fa31b466bb473797f0d0314c0bdf, 168'h00e2977c479e6d25703cebbc6bd561938cc9d1bfb9},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=168b(21B), s=168b(21B)
  '{375, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h4cbacc728670e4e1df367749fce32c6a4f17bc634bc52f502d44cc95, 232'h00e0a864b52cdffddaeb70ed9f073484a45858889c58e80ec8007e9fc6, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{376, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h4cbacc728670e4e1df367749fce32c6a4f17bc634bc52f502d44cc95, 232'h00e0a864b52cdffddaeb70ed9f073484a45858889c58e80ec8007e9fc6, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 8'h00},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{377, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h4b9c0cf9f218f64d1317ffc18caf11797cbb431550816b42e658da6c, 224'h5051333576ab8be2753bcfbad797b29c0b8eb76b4b310bb24f3c6ec7, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h74d89d2b42107a17e0df7430a84102f0c3befe18e59ea9ed5aef3195},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{378, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008981be0db57c743232f8a5d30b419840c4d38087d66c501597f737ac, 232'h00b07a341cac19c626da4adb9f3119cb4439e954b1718a7eae45f7a933, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h2a179e7ed670727c33ba8da63fe226140a7fcf62d2cfaea7ea59d1d4},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{379, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h69f46cfddcec6520e4e65590c64466c19cff0f581e13ed401d4f3470, 232'h00cfb829ac4e52055461d0785876d78e3d5889a7749be663a6bf08459b, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h6d50b1cb505189520a6901a895ea13458ff5076156c27efc00639c35},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{380, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0086ae72267749417993992aa8724e9d760dc3962b2ad01ebc28019fa0, 224'h5a107cf5332ff42f5516451f2298a362a894d95ba849d48ed389ffd5, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h0f59ae2e4259dbe0997caabcdb25bdbe8d6df67f433a4651342d5219},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{381, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d39979285ed39d2250c5125305868dbd4274b8a603d571e3537c2ea5, 232'h00f7c67e822535efc4c1021b6b312c34e4d60be2e89984e95f5dddb7de, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h5e10dd8d9f91876988f21a2bc2fefa4df57ab4efc82ca41a773ae802},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{382, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h5329099622fe9e1008c891fff3ba768c6d764d420509fd232830603b, 224'h2d9d32aff3af504eb4389dc7bde4f9c4c5fdac7bff001d6da369104c, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h511eb0edc14410a1c38d655e04e0c99cd8af84d8caa0ffd69da2dc44},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{383, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0090d1161f4794186cc6d0baeaa03f63e84ae61b3428712cd561978ecd, 232'h00acd7e006ada0004b6ea0f27da9ea26791a94292e57e3584af0de87c5, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h11577274428aaa4ac5d23552e64d35c2e45667773fe77fba629f873f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{384, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h326aa12c68fd569b573884a97b899c197c18fb9c509782be8b18011f, 232'h0082d76e993348dd4de2440a6d7bbfcd7461729a6ac70a3fade02fbd8b, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h2fb159d4c8769a346ee620bb1e5027f2aa0fd3b1d8b3a2411c9b9ca0},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{385, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h0633d37de65ad8897f863b485babc75cb14175692597db295e4d2beb, 224'h649f25584f8f9f3121549431e1e3ea5290ed186d443ac4b53df57b14, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h59d3622af6be99859f0aea85aa20e669ec373992af2856f37dea777f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{386, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0093f80c5d235dbb8efb8622bf70716316b021ece8a37d2ff33a422cbd, 232'h00b0fe70e8e87e04736a54a943d524b3ef27628d7f7688e901fdb25f40, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h3296bcaf337a66617b38e2ab65833612cd0bae1b7b3e670863dac215},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{387, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h6bd84040f3c08088a7dab45cb4a455a8b5336a00f2b2899779adc048, 232'h00cf5d1bdbb1042789adeb363dbd7c4f776560f7d3c6ff24e58d0709c0, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h1b468ea6fa697becc552ec879c3e9ffdd72969403d5fb745bbd7f366},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{388, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h6a942adc74e5a542beb5a9ed73166bba16a621fde05fad8feb93041a, 232'h00b9d8e5797a2e237b2785c36f24156dd40d3ed35064f8878bb6db114a, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h244b2ee0f3acf3ca0d086215fbc12728516ffc93c03d27a601d31a8a},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{389, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h74897882013164324092db05bb1d2e0d44386fea0ad1b2eefec19565, 224'h0f28f541785399eb1b825131e82b18da9a30049686fd4af36fff43ce, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h5625c3f523582b7986ad997a8488acfbfc4b2db75913a1fa4b437ec5},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{390, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0081a4a2c2c959ba5ef743d32f173b1e24567ea1c37fc5cf6e36b02577, 224'h079d37fa3c2f8540bed4d6465ff45ed71878ba86cee8ffb4776231ad, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b55, 224'h148bd1fd5c6502009ef1febb26c374cacd3a62e7f3f232e21f145115},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{396, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c73ef8ec74b35b83942ec13f90b838147e31e00c84c82166fbee4a8e, 224'h2adf5032da443a8ec22a4cff4c3a4724a79ace6394048237b5bd6890, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b4e, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b4e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{399, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h14d87a664bac68655b1767aec2bb50c920f92c31eb07d4f08cefd2b2, 224'h618d1fbfff7dfa24e85b3ac5de8e433618fe56480698113a76915f80, 40'h0100001a90, 224'h050bc5eda83286e4e8506020be6a8eb2d500ea3be9104339e91396fc},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{404, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d67cb3bb26f994c8a6e591b821245f5e118b2667b7f75c9251eef200, 224'h61b5696a63106e89fd531b9ccdfae032a668fe274bc1cbf5be1bc200, 40'h0100001a90, 224'h12b14ca9894b5a17a0c6db3c25795ee7825cdea7d37ffcbbcc8b03df},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{406, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h04f39a7ded5b62d429e3af6d2718457ffd87a9d00f4b5389e0230848, 224'h57b0cbadb8326c12a2fc15a42206d515011ec6e5272583e5d2036c1e, 40'h0100001a90, 224'h2dc3c8b28aecf3beb728695c47ea27593723a6811531134649fd0ffb},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=40b(5B), s=224b(28B)
  '{409, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a824ae928cb209d3d4143a8cd10a7b29d863150a5482f873972e6031, 224'h12f9d12f2fff94f4e0a5b9e3e5a88bc21b2d09da15584ca655c31094, 40'h0100001a90, 32'h55555e30},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=40b(5B), s=32b(4B)
  '{411, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h5e423679db282576cec351f1500a4ee1a3e6bc146b76c147c3798fe3, 232'h00ed029bdb0474eddaad50e2a6f2780ff184b33f4c38c03738ed6c1ba7, 40'h0100001a90, 224'h39232f26cb0fcd6b2eeb69ba41b9ef00813616da98cd16e2ef21123f},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=40b(5B), s=224b(28B)
  '{412, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h038925a04a7e62c3f709ae4150051692290405fc3e2c0ec2eb0de428, 232'h008d7148d65237c36fe18e125447adf9189793b86f5256e915c52d44d9, 40'h0100001a90, 224'h121c0384a8d015f000000000000021bc8ed98db7f846a8b77b820ac0},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=40b(5B), s=224b(28B)
  '{422, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h5126d8509cc88bd0ae29c97062b8ba4b416906294a9331bc678dd362, 224'h65171023f5de2d1c8a2da0080f50b29972875fc7c1bf9428d95aa704, 224'h5555555555555555555555555555f44d9ba4208198fae325d2353b52, 224'h33333333333333333333333333339294f6fc1380f5635516b1532397}  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224K1_SHA256_V1_SV
