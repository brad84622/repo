`ifndef WYCHERPROOF_SECP224R1_SHA224_SV
`define WYCHERPROOF_SECP224R1_SHA224_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224r1_sha224;

localparam int TEST_VECTORS_SECP224R1_SHA224_NUM = 60;

ecdsa_vector_secp224r1_sha224 test_vectors_secp224r1_sha224 [] = '{
  '{1, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'h2840bf24f6f66be287066b7cbf38788e1b7770b18fd1aa6a26d7c6dc},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{2, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'hd7bf40db0909941d78f9948340c69e14c5417f8c840b7edb35846361},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{115, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 0},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=0b(0B)
  '{124, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'h00d7bf40db0909941d78f9948340c69e14c5417f8c840b7edb358463},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{130, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{139, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'hd7bf40db0909941d78f9948340c78771e4888f4e702e5595d9283924},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{143, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h70049af31f8348673d56cece2b27e587a402f2a48f0b21a7911a480a, 224'h2840bf24f6f66be287066b7cbf3961eb3abe80737bf48124ca7b9c9f},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{144, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{230, 1'b1, 224'h45dbc3e1ba272f7770c91d10827c5b55efd21f769e8c16c22d50d4da, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h326bc06353f7f9c9f77b8f4b55464e8619944e7879402cca572e041a, 224'h3116e1a38e4ab2008eca032fb2d185e5c21a232eaf4507ae56177fd2},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{235, 1'b1, 224'h75a5fb77bbf26e1d0000000032c79994621210a6548b17196169f7a6, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h2b98c67ebf6597b08bc7f1b73ff8662cf125e9700ec973ece9c6ff48, 224'h2e3f72a8f76e12c8cdf4487e0956c1ef4578e1da4d29d8db824d415b},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{240, 1'b1, 224'h4bb4c6ef041cc67b6d219b8bb8efde000000004ed8c91a45116088a1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h64c084f6b775bbf7915c1964a68b0259629328598f13557872867830, 224'h2a6f3b289d130ec3d99e4caaf601497895a069c1a5a75b559ad28444},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{245, 1'b1, 224'h164913b0ffffffff8271b08e9f2f12b2d2f280c4bcfa2e10cf3bcdef, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5dfc6fad385bdb24b2b70a64fd4253405c0028bb36f4793aa3bd31fe, 224'h1c210b74924171378992b03bb1bd78c5cfcfc879d2e5c736d35516c3},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{247, 1'b1, 224'ha6f97a37213effffffff1ee90d31e0879292f54edb4ecd18a8de16f1, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h120055f90ad1290c4c5fc5faf69b215139182c770d2b55e95712442f, 224'h01ac47f7446543d4003b039d9f54daa9d0799f98291a32df4fcd472a},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{249, 1'b1, 224'ha547b8919fb96574b64e1689ffffffff92bc14d17ee24df64421cf21, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h57daddb0cb6af939b1ea1aaf4bc72e56150c0c46a581827193e65d17, 224'h3bc37bde4e60b789ba86a054d37f1191e0814926c1a0100168d16c17},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{250, 1'b1, 224'h51a094b7010ba80e7b697b1455ffffffff5eec554b8f0fbca92e6384, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3a74102bd1fc617018efc4fbc042e719a81b55830aac1f1dcdedec65, 224'h4bb9fe90015a45f31c8c95dda24f54fcdb64682c13f68d4da3d1abe0},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{252, 1'b1, 224'h324c363aa6df32aded1b26d162c72bcaffffffff00b71dc4e28f991e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3c212b5a7e65d9af44643bd62fa42a9b9cffe6bdb623e9b9e4337156, 224'h29c8121a12427a324e5d551ff5a83d3c252e32257af2800d080817d2},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{253, 1'b1, 224'hfe1211e72fe25ef2f8b531b268553f6835b5ffffffff72b5d98c3d83, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1630554989fffd0e35f2d9105623d73a543634c48000484c422272ca, 224'h214da487d5e51f73814dff80a08c77bd8a83a9889a1b26a5578ba954},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{260, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00ea3ea2873b6fc099bfd779b0a2c23c2c4354e2fec4536f3b8e420988, 232'h00f97e1c7646b4eb3de616752f415ab3a6f696d1d674fb4b6732252382, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{262, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00b157315cc1aaeae64eb5b38452884195fdfe8a15fb5618284f48afe5, 232'h00e1fbbaad729477a45f3752b7f72ad2f9cd7dce4158a8e21b8127e8a7, 8'h03, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{263, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h0087d9d964044b5b16801f32de9f3f9066194e8bf80affa3cb0d4ddb1d, 232'h00b5eb9b6594e6d1bcacd0fd9d67c408f789dfb95feb79a6e2fb9c4cee, 8'h03, 8'h03},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{264, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h461b435af09ede35e74dac21f9af7b1b9998213039f8785d4a4905f5, 224'h18b89bde69de34a482638461d09386e7193ca90ca5b3038e2a3885d1, 8'h03, 8'h04},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{268, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00beb9d8dcba48146b9032688ecea947a231e7d0e6ce17d76b56ed6348, 224'h35503f3b4af414870ef03383784b1d846b3e07b8e9fc2d6190a3bfda, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{269, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h1955ba3f90e7a739471a5d182b594c9747eb49d5356203f3bb8b939c, 232'h00807d88ce3a0885bfa5b5b7f6e9beb18285e7130524b6c1498b3269ee, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{273, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00b671296dd5f690502e4b1500e4acb4c82d3aa8dfbc5868a643f86a3c, 232'h00a46ba8c3a7b823259522291e2416232276cca8503cc8dbf941f1d93d, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{274, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00b671296dd5f690502e4b1500e4acb4c82d3aa8dfbc5868a643f86a3c, 232'h00a46ba8c3a7b823259522291e2416232276cca8503cc8dbf941f1d93d, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{275, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h76e34b57a8c61df59cb0b7921cec6e5422344033f7accb7b3179e682, 232'h00cefd0a848309d1decf98a3b9e333691b95c17821cb681137630c02e2, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{276, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h51839e545c872f4a381f278ed5b4c24cf38aac77b02953405618bf27, 224'h394e41226594c499db6a7dd7a6901bda5e6474b1ffa10a6567210010, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{277, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00a3ec90053d1e100815d1becfe96c9b3646e52df794f6b03b766a7574, 232'h00c3b7e17e73acc8cefe71b6eb13d4f1c94c57e58bee43c69d9d41a964, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{278, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00b5c09b4851a67371eee7bbf02451e5208c40de61bc1a33df2710b384, 232'h00dcce4e5b83c32a800e8de28fa936d582cdcad185e894caac797f1d14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{280, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h43c9ccd08a80bca18022722b0bdcd790d82a3ef8b65c3f34204bb472, 232'h009ee1c1f00598130b2313a3e38a3798d03dac665cff20f36ce8a2024a, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{283, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h3d2e9bb9a712bf3ad42ac30659fdbda9be9956537f9f37cd05f0ff37, 224'h7d5982d6d9266d774942c44d9eb3501051d3b9688610131e7856ef36, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7ac54a381d9bd3f2698359d6f658b5e4167d15a75b576e82d2efbd37},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{284, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00a0be2f10144b9b42b016f1bd9fca30e4c24aae4775596c7cdb07ae60, 232'h00d60ff3a70f1541631f6087d3f3b3fe376d2305b50b94821106412479, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h4fbb063e82402e16fe14edda4d7986b0b88344a1f53b0e2684ee7e31},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{290, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h3c59e13982fd9c1a45991b1e9d79e939a52a62ca479764f1477e2813, 224'h1b004c9bffd7f00c05e3168c625cc93ab7a0f1ba8d6fa26a4d5162cb, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2e416eaa8279952a0d6ba4eb13cbfee69cf7bcae437232fbfa5a5d5b},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{293, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h4108e0ccd47cba09fb7ed4d9f3455823780965157861c1bf8f93d34b, 224'h46d6fdb71e9e89adaae71376b13fd17644b11eed00d498783da0ba1a, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{295, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h7dc09710f4f586af05b08f0c9dcd48b1308733c97767fc286d1c7283, 224'h4353a704c7950b8f4a11394bc8db06adccf19d8ed95c7f214a173137, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{297, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00e012dc20cca5bd2adfaa27f57419596ce09ed0f18a9148e30a0f6ed2, 224'h55beca1b5e3e2485ef9537ae48a67b72dbcf6d7b33372023a5c443e8, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{299, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h08a6e167536a47aaa224fec21ce077642efdb97d93ae16b9672279f4, 224'h33fb9f1abb25f2c0c3e6008ac857ede4a89ca8d9d08b8996614969ac, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{301, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h2d59efd841a44b83fd42e6a2984a53fa93ad242c11678f92202cccfb, 232'h0095bcaf0b2f6eb0e6d4d83e3260e037d3dc0e48ab6c4141ce6b56cad0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{302, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h1161c7add6f67f995b93e19eb18bd5e73fd71d6bb10dceef0b792e9c, 224'h08c44cef9826b4ed67508c09d07ec857a0ea49ed1a7f1fa2c74cb838, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{306, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00e2ef8c8ccb58eba287d9279b349e7652cca3e7cda188a5f179d77142, 232'h00f87594f3664c0faf7b59670e353a370d1d68ad89d6a1e246b4d03bee, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{307, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00b8bf3ef9646abfffb84220104ec996a92cef33f9328ec4cb1ea69948, 224'h4fea51a0de9e9d801babd42ca0924b36498bc5900fbeb9cbd5ad9c1a, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{309, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h5599a3faf96aba7302bd3d98cfde69525b7292762383f4a0b5c31039, 224'h3faa45feb6c35d2b7bf25ffc633c420ebfc4e715765302c5a11ac793, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{311, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00aced4ea8949e5ae37ef2f5eb5e00675d08e17c34be6677b0f269b672, 224'h5e3ad0af49ebfff415ee4f2a838ead1f84cafaa652c17acc26130725, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{312, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h3e8c1bcc16195e8769e25d4c859807dffe178bed5bca9db06efa1532, 224'h4e3b53b3048b8ccd8cdc1265be240c8ee204060486a99ad31eaad3a4, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=224b(28B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{319, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=224b(28B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{321, 1'b0, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{325, 1'b1, 224'h753bb40078934081d7bd113ec49b19ef09d1ba33498690516d4d122c, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h01ec1ff15c8a55d697a5424d674753f82f711593828368d2fbb41a17, 224'h20d9089db7baf46b8135e17e01645e732d22d5adb20e3772da740eee},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 224'hbd4f57a4cfb1649cca33372f5c5ad32b993ff73aaf4fb75d52798480, 224'h4c246670658a1d41f5d77bce246cbe386ac22848e269b9d4cd67c466, 232'h00ddd947153d39b2d42533a460def26880408caf2dd3dd48fe888cd176, 224'h3e46e9ba4dc089ff30fa8c0209c31b11ff49dbeec090f9f53c000c75, 224'h6f2e3b36369416602bca83206809ed898fcf158a56c25a5474143f68},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{338, 1'b1, 224'h3dc6a3fd912b08bf15170296c4f1694f512ffa1dc9bddb8b9e1c8d38, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h576bb86c517bfecdc930a4c8501725548d425afbb96d93f5c1e2a0e1, 224'h77248c5ecd620c431438c50e6bee6858091b54a87f8548ae35c21027},  // lens: hash=224b(28B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 224'h3dc6a3fd912b08bf15170296c4f1694f512ffa1dc9bddb8b9e1c8d38, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 192'h762d28f1fdc219184f81681fbff566d465b5f1f31e872df5, 224'h2558a42e79689244bccd5e855f6a1e42b4ff726873f30b532b89ef53, 224'h07f9bd947785187175d848b6e2d79f7ab3bbc1087b42590b0cfb256a},  // lens: hash=224b(28B), x=224b(28B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{344, 1'b1, 224'h3dc6a3fd912b08bf15170296c4f1694f512ffa1dc9bddb8b9e1c8d38, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h305ccf0b5d0cf33dc745bb7c7964c233f6cfd8892a1c1ae9f50b2f3f, 224'h785f6e85f5e652587c6e15d0c45c427278cf65bb1429a57d8826ca39},  // lens: hash=224b(28B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{347, 1'b1, 224'h3dc6a3fd912b08bf15170296c4f1694f512ffa1dc9bddb8b9e1c8d38, 200'h00f7e4713d085112112c37cdf4601ff688da796016b71a727a, 232'h00de5a9ec165054cc987f9dc87e9991b92e4fa649ca655eeae9f2a30e1, 224'h0e05ed675c673e5e70a4fdd5a47b114c5d542d4f6d7a367597d713ea, 224'h26d70d65c48430373363987810bdcc556e02718eab214403ae008db4}  // lens: hash=224b(28B), x=200b(25B), y=232b(29B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224R1_SHA224_SV
