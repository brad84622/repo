`ifndef WYCHERPROOF_SECP256K1_SHA256_P1363_SV
`define WYCHERPROOF_SECP256K1_SHA256_P1363_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp256k1_sha256_p1363;

localparam int TEST_VECTORS_SECP256K1_SHA256_P1363_NUM = 207;

ecdsa_vector_secp256k1_sha256_p1363 test_vectors_secp256k1_sha256_p1363 [] = '{
  '{1, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h813ef79ccefa9a56f7ba805f0e478584fe5f0dd5f567bc09b5123ccbc9832365, 256'h900e75ad233fcc908509dbff5922647db37c21f4afd3203ae8dc4ae7794b0f87},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{3, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7ec10863310565a908457fa0f1b87a79bc4fcf10b9e0e4320ac021c106b31ddc, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{5, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h7ec10863310565a908457fa0f1b87a7b01a0f22a0a9843f64aedc334367cdc9b, 256'h6ff18a52dcc0336f7af62400a6dd9b810732baf1ff758000d6f613a556eb31ba},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{8, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h813ef79ccefa9a56f7ba805f0e478584fe5f0dd5f567bc09b5123ccbc9832365, 256'h900e75ad233fcc908509dbff5922647ef8cd450e008a7fff2909ec5aa914ce46},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{9, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{10, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{11, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{12, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{13, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{14, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{15, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000000, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{16, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{17, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{18, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{19, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{20, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{21, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{22, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{23, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{24, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{25, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{26, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{27, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{28, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{29, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{30, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{31, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{32, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{33, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{34, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{35, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{36, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{37, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{38, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{39, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{40, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{41, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{42, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{43, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{44, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{45, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{46, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{47, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{48, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{49, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{50, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{51, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{52, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{53, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364141},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{54, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364140},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{55, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{56, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{57, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc30},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{58, 1'b1, 256'hb78f33ca6d031315ab4c29b4429e6e8f8978517d49192c90fb2266bea6842918, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hdd1b7d09a7bd8218961034a39a87fecf5314f00c4d25eb58a07ac85e85eab516, 256'h35138c401ef8d3493d65c9002fe62b43aee568731b744548358996d9cc427e06},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{59, 1'b1, 256'h00000000690ed426ccf17803ebe2bd0884bcd58a1bb5e7477ead3645f356e7a9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h95c29267d972a043d955224546222bba343fc1d4db0fec262a33ac61305696ae, 256'h6edfe96713aed56f8a28a6653f57e0b829712e5eddc67f34682b24f0676b2640},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{60, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h28f94a894e92024699e345fe66971e3edcd050023386135ab3939d550898fb25, 256'hcd69c1a42be05a6ee1270c821479251e134c21858d800bda6f4e98b37196238e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{61, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hbe26b18f9549f89f411a9b52536b15aa270b84548d0e859a1952a27af1a77ac6, 256'h8f3e2b05632fc33715572af9124681113f2b84325b80154c044a544dc1a8fa12},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{62, 1'b1, 256'h67ab1900000000784769c4ecb9e164d6642b8499588b89855be1ec355d0841a0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hb1a4b1478e65cc3eafdf225d1298b43f2da19e4bcff7eacc0a2e98cd4b74b114, 256'he8655ce1cfb33ebd30af8ce8e8ae4d6f7b50cd3e22af51bf69e0a2851760d52b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{63, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h325332021261f1bd18f2712aa1e2252da23796da8a4b1ff6ea18cafec7e171f2, 256'h40b4f5e287ee61fc3c804186982360891eaa35c75f05a43ecd48b35d984a6648},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{64, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'ha23ad18d8fc66d81af0903890cbd453a554cb04cdc1a8ca7f7f78e5367ed88a0, 256'hdc1c14d31e3fb158b73c764268c8b55579734a7e2a2c9b5ee5d9d0144ef652eb},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{65, 1'b1, 256'h9b6cd3b812610000000026941a0f0bb53255ea4c9fd0cb3426e3a54b9fc6965c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2bdea41cda63a2d14bf47353bd20880a690901de7cd6e3cc6d8ed5ba0cdb1091, 256'hc31599433036064073835b1e3eba8335a650c8fd786f94fe235ad7d41dc94c7a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{66, 1'b1, 256'h883ae39f50bf0100000000e7561c26fc82a52baa51c71ca877162f93c4ae0186, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hd7cd76ec01c1b1079eba9e2aa2a397243c4758c98a1ba0b7404a340b9b00ced6, 256'hca8affe1e626dd192174c2937b15bc48f77b5bdfe01f073a8aeaf7f24dc6c85b},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{67, 1'b1, 256'ha1ce5d6e5ecaf28b0000000000fa7cd010540f420fb4ff7401fe9fce011d0ba6, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'ha872c744d936db21a10c361dd5c9063355f84902219652f6fc56dc95a7139d96, 256'h400df7575d9756210e9ccc77162c6b593c7746cfb48ac263c42750b421ef4bb9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{68, 1'b1, 256'h8ea5f645f373f580930000000038345397330012a8ee836c5494cdffd5ee8054, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h9fa9afe07752da10b36d3afcd0fe44bfc40244d75203599cf8f5047fa3453854, 256'haf1f583fec4040ae7e68c968d2bb4b494eec3a33edc7c0ccf95f7f75bc2569c7},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{69, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h885640384d0d910efb177b46be6c3dc5cac81f0b88c3190bb6b5f99c2641f205, 256'h738ed9bff116306d9caa0f8fc608be243e0b567779d8dab03e8e19d553f1dc8e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{70, 1'b1, 256'hd0462673154cce587dde8800000000e98d35f1f45cf9c3bf46ada2de4c568c34, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2d051f91c5a9d440c5676985710483bc4f1a6c611b10c95a2ff0363d90c2a458, 256'h92206b19045a41a797cc2f3ac30de9518165e96d5b86341ecb3bcff231b3fd65},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{71, 1'b1, 256'hbd90640269a7822680cedfef000000000caef15a6171059ab83e7b4418d7278f, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hf3ac2523967482f53d508522712d583f4379cd824101ff635ea0935117baa54f, 256'h27f10812227397e02cea96fb0e680761636dab2b080d1fc5d11685cbe8500cfe},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{72, 1'b1, 256'h33239a52d72f1311512e41222a00000000d2dcceb301c54b4beae8e284788a73, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h96447cf68c3ab7266ed7447de3ac52fed7cc08cbdfea391c18a9b8ab370bc913, 256'hf0a1878b2c53f16e70fe377a5e9c6e86f18ae480a22bb499f5b32e7109c07385},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{73, 1'b1, 256'hb8d64fbcd4a1c10f1365d4e6d95c000000007ee4a21a1cbe1dc84c2d941ffaf1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h530a0832b691da0b5619a0b11de6877f3c0971baaa68ed122758c29caaf46b72, 256'h93761bb0a14ccf9f15b4b9ce73c6ec700bd015b8cb1cfac56837f4463f53074e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{74, 1'b1, 256'h01603d3982bf77d7a3fef3183ed092000000003a227420db4088b20fe0e9d84a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h9c54c25500bde0b92d72d6ec483dc2482f3654294ca74de796b681255ed58a77, 256'h988bac394a90ad89ce360984c0c149dcbd2684bb64498ace90bcf6b6af1c170e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{75, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'he7909d41439e2f6af29136c7348ca2641a2b070d5b64f91ea9da7070c7a2618b, 256'h42d782f132fa1d36c2c88ba27c3d678d80184a5d1eccac7501f0b47e3d205008},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{76, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5924873209593135a4c3da7bb381227f8a4b6aa9f34fe5bb7f8fbc131a039ffe, 256'he0e44ee4bbe370155bf0bbdec265bf9fe31c0746faab446de62e3631eacd111f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{77, 1'b1, 256'h307bfaaffb650c889c84bf83f0300e5dc87e000000008408fd5f64b582e3bb14, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'heeb692c9b262969b231c38b5a7f60649e0c875cd64df88f33aa571fa3d29ab0e, 256'h218b3a1eb06379c2c18cf51b06430786d1c64cd2d24c9b232b23e5bac7989acd},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{78, 1'b1, 256'hbab5c4f4df540d7b33324d36bb0c157551527c00000000e4af574bb4d54ea6b8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'ha40034177f36091c2b653684a0e3eb5d4bff18e4d09f664c2800e7cafda1daf8, 256'h3a3ec29853704e52031c58927a800a968353adc3d973beba9172cbbeab4dd149},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{79, 1'b1, 256'hd4ba47f6ae28f274e4f58d8036f9c36ec2456f5b00000000c3b869197ef5e15e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hb5d795cc75cea5c434fa4185180cd6bd21223f3d5a86da6670d71d95680dadbf, 256'hab1b277ef5ffe134460835e3d1402461ba104cb50b16f397fdc7a9abfefef280},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{80, 1'b1, 256'h79fd19c7235ea212f29f1fa00984342afe0f10aafd00000000801e47f8c184e1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h07dc2478d43c1232a4595608c64426c35510051a631ae6a5a6eb1161e57e42e1, 256'h4a59ea0fdb72d12165cea3bf1ca86ba97517bd188db3dbd21a5a157850021984},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{81, 1'b1, 256'h8c291e8eeaa45adbaf9aba5c0583462d79cbeb7ac97300000000a37ea6700cda, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hddd20c4a05596ca868b558839fce9f6511ddd83d1ccb53f82e5269d559a01552, 256'ha46e8cb8d626cf6c00ddedc3b5da7e613ac376445ee260743f06f79054c7d42a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{82, 1'b1, 256'h0eaae8641084fa979803efbfb8140732f4cdcf66c3f78a000000003c278a6b21, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h9cde6e0ede0a003f02fda0a01b59facfe5dec063318f279ce2de7a9b1062f7b7, 256'h2886a5b8c679bdf8224c66f908fd6205492cb70b0068d46ae4f33a4149b12a52},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{83, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hc5771016d0dd6357143c89f684cd740423502554c0c59aa8c99584f1ff38f609, 256'hab4bfa0bb88ab99791b9b3ab9c4b02bd2a57ae8dde50b9064063fcf85315cfe5},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{84, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'ha24ebc0ec224bd67ae397cbe6fa37b3125adbd34891abe2d7c7356921916dfe6, 256'h34f6eb6374731bbbafc4924fb8b0bdcdda49456d724cdae6178d87014cb53d8c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{85, 1'b1, 256'h62aac98818b3b84a2c214f0d5e72ef286e1030cb53d9a82b690e00000000cd15, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2557d64a7aee2e0931c012e4fea1cd3a2c334edae68cdeb7158caf21b68e5a24, 256'h80f93244956ffdc568c77d12684f7f004fa92da7e60ae94a1b98c422e23eda34},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{86, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hc4f2eccbb6a24350c8466450b9d61b207ee359e037b3dcedb42a3f2e6dd6aeb5, 256'hcd9c394a65d0aa322e391eb76b2a1a687f8620a88adef3a01eb8e4fb05b6477a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{87, 1'b1, 256'h0da0a1d2851d33023834f2098c0880096b4320bea836cd9cbb6ff6c800000000, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'heff04781c9cbcd162d0a25a6e2ebcca43506c523385cb515d49ea38a1b12fcad, 256'hea5328ce6b36e56ab87acb0dcfea498bcec1bba86a065268f6eff3c41c4b0c9c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{88, 1'b1, 256'hffffffff293886d3086fd567aafd598f0fe975f735887194a764a231e82d289a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hf58b4e3110a64bf1b5db97639ee0e5a9c8dfa49dc59b679891f520fdf0584c87, 256'hd32701ae777511624c1f8abbf02b248b04e7a9eb27938f524f3e8828ba40164a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{89, 1'b1, 256'h7bffffffff2376d1e3c03445a072e24326acdc4ce127ec2e0e8d9ca99527e7b7, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hf8abecaa4f0c502de4bf5903d48417f786bf92e8ad72fec0bd7fcb7800c0bbe3, 256'h4c7f9e231076a30b7ae36b0cebe69ccef1cd194f7cce93a5588fd6814f437c0e},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{90, 1'b1, 256'ha2b5ffffffffebb251b085377605a224bc80872602a6e467fd016807e97fa395, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5d5b38bd37ad498b2227a633268a8cca879a5c7c94a4e416bd0a614d09e606d2, 256'h12b8d664ea9991062ecbb834e58400e25c46007af84f6007d7f1685443269afe},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{91, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0c1cd9fe4034f086a2b52d65b9d3834d72aebe7f33dfe8f976da82648177d8e3, 256'h13105782e3d0cfe85c2778dec1a848b27ac0ae071aa6da341a9553a946b41e59},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{92, 1'b1, 256'h958415d8ffffffffabad03e2fc662dc3ba203521177502298df56f36600e0f8b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hae7935fb96ff246b7b5d5662870d1ba587b03d6e1360baf47988b5c02ccc1a5b, 256'h5f00c323272083782d4a59f2dfd65e49de0693627016900ef7e61428056664b3},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{93, 1'b1, 256'hf1d8de4858ffffffff1281093536f47fe13deb04e1fbe8fb954521b6975420f8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h00a134b5c6ccbcefd4c882b945baeb4933444172795fa6796aae149067547098, 256'ha991b9efa2db276feae1c115c140770901839d87e60e7ec45a2b81cf3b437be6},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{94, 1'b1, 256'h0927895f2802ffffffff10782dd14a3b32dc5d47c05ef6f1876b95c81fc31def, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2e4721363ad3992c139e5a1c26395d2c2d777824aa24fde075e0d7381171309d, 256'h8bf083b6bbe71ecff22baed087d5a77eaeaf726bf14ace2c03fd6e37ba6c26f2},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{95, 1'b1, 256'h60907984aa7e8effffffff4f332862a10a57c3063fb5a30624cf6a0c3ac80589, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h6852e9d3cd9fe373c2d504877967d365ab1456707b6817a042864694e1960ccf, 256'hf9b4d815ebd4cf77847b37952334d05b2045cb398d4c21ba207922a7a4714d84},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{96, 1'b1, 256'hc6ff198484939170ffffffff0af42cda50f9a5f50636ea6942d6b9b8cd6ae1e2, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h188a8c5648dc79eace158cf886c62b5468f05fd95f03a7635c5b4c31f09af4c5, 256'h36361a0b571a00c6cd5e686ccbfcfa703c4f97e48938346d0c103fdc76dc5867},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{97, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'ha74f1fb9a8263f62fc4416a5b7d584f4206f3996bb91f6fc8e73b9e92bad0e13, 256'h6815032e8c7d76c3ab06a86f33249ce9940148cb36d1f417c2e992e801afa3fa},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{98, 1'b1, 256'h6f0e3eeaf42b28132b88fffffffff6c8665604d34acb19037e1ab78caaaac6ff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h07244865b72ff37e62e3146f0dc14682badd7197799135f0b00ade7671742bfe, 256'hf27f3ddc7124b1b58579573a835650e7a8bad5eeb96e9da215cd7bf9a2a039ed},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{99, 1'b1, 256'hcdb549f773b3e62b3708d1ffffffffbe48f7c0591ddcae7d2cb222d1f8017ab9, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hda7fdd05b5badabd619d805c4ee7d9a84f84ddd5cf9c5bf4d4338140d689ef08, 256'h28f1cf4fa1c3c5862cfa149c0013cf5fe6cf5076cae000511063e7de25bb38e5},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{100, 1'b1, 256'h2c3f26f96a3ac0051df4989bffffffff9fd64886c1dc4f9924d8fd6f0edb0484, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hd3027c656f6d4fdfd8ede22093e3c303b0133c340d615e7756f6253aea927238, 256'hf6510f9f371b31068d68bfeeaa720eb9bbdc8040145fcf88d4e0b58de0777d2a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{101, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0bf6c0188dc9571cd0e21eecac5fbb19d2434988e9cc10244593ef3a98099f69, 256'h4864a562661f9221ec88e3dd0bc2f6e27ac128c30cc1a80f79ec670a22b042ee},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{102, 1'b1, 256'h4f9618f98e2d3a15b24094f72bb5ffffffffa2fd3e2893683e5a6ab8cf0ee610, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'hae459640d5d1179be47a47fa538e16d94ddea5585e7a244804a51742c686443a, 256'h6c8e30e530a634fae80b3ceb062978b39edbe19777e0a24553b68886181fd897},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{103, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h1cf3517ba3bf2ab8b9ead4ebb6e866cb88a1deacb6a785d3b63b483ca02ac495, 256'h249a798b73606f55f5f1c70de67cb1a0cff95d7dc50b3a617df861bad3c6b1c9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{104, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'he69b5238265ea35d77e4dd172288d8cea19810a10292617d5976519dc5757cb8, 256'h4b03c5bc47e826bdb27328abd38d3056d77476b2130f3df6ec4891af08ba1e29},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{105, 1'b1, 256'h3c80de54cd9226989443d593fa4fd6597e280ebeffffffffc1847eb76c217a95, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5f9d7d7c870d085fc1d49fff69e4a275812800d2cf8973e7325866cb40fa2b6f, 256'h6d1f5491d9f717a597a15fd540406486d76a44697b3f0d9d6dcef6669f8a0a56},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{106, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h0a7d5b1959f71df9f817146ee49bd5c89b431e7993e2fdecab6858957da685ae, 256'h0f8aad2d254690bdc13f34a4fec44a02fd745a422df05ccbb54635a8b86b9609},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{107, 1'b1, 256'h8f65d92927cfb86a84dd59623fb531bb599e4d5f7289ffffffff2f1f2f57881c, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h79e88bf576b74bc07ca142395fda28f03d3d5e640b0b4ff0752c6d94cd553408, 256'h32cea05bd2d706c8f6036a507e2ab7766004f0904e2e5c5862749c0073245d6a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{108, 1'b1, 256'h6b63e9a74e092120160bea3877dace8a2cc7cd0e8426cbfffffffffafc8c3ca8, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h9d54e037a00212b377bc8874798b8da080564bbdf7e07591b861285809d01488, 256'h18b4e557667a82bd95965f0706f81a29243fbdd86968a7ebeb43069db3b18c7f},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{109, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h2664f1ffa982fedbcc7cab1b8bc6e2cb420218d2a6077ad08e591ba9feab33bd, 256'h49f5c7cb515e83872a3d41b4cdb85f242ad9d61a5bfc01debfbb52c6c84ba728},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{110, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h5827518344844fd6a7de73cbb0a6befdea7b13d2dee4475317f0f18ffc81524b, 256'hb0a334b1f4b774a5a289f553224d286d239ef8a90929ed2d91423e024eb7fa66},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{111, 1'b1, 256'h08fb565610a79baa0c566c66228d81814f8c53a15b96e602fb49ffffffffff6e, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h97ab19bd139cac319325869218b1bce111875d63fb12098a04b0cd59b6fdd3a3, 256'hbce26315c5dbc7b8cfc31425a9b89bccea7aa9477d711a4d377f833dcc28f820},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{112, 1'b1, 256'hd59291cc2cf89f3087715fcb1aa4e79aa2403f748e97d7cd28ecaefeffffffff, 264'h00b838ff44e5bc177bf21189d0766082fc9d843226887fc9760371100b7ee20a6f, 264'h00f0c9d75bfba7b31a6bca1974496eeb56de357071955d83c4b1badaa0b21832e9, 256'h52c683144e44119ae2013749d4964ef67509278f6d38ba869adcfa69970e123d, 256'h3479910167408f45bda420a626ec9c4ec711c1274be092198b4187c018b562ca},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{113, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h07310f90a9eae149a08402f54194a0f7b4ac427bf8d9bd6c7681071dc47dc362, 256'h26a6d37ac46d61fd600c0bf1bff87689ed117dda6b0e59318ae010a197a26ca0, 256'h000000000000000000000000000000014551231950b75fc4402da1722fc9baeb, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{114, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h07310f90a9eae149a08402f54194a0f7b4ac427bf8d9bd6c7681071dc47dc362, 256'h26a6d37ac46d61fd600c0bf1bff87689ed117dda6b0e59318ae010a197a26ca0, 256'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffefffffc2c, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{115, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00bc97e7585eecad48e16683bc4091708e1a930c683fc47001d4b383594f2c4e22, 256'h705989cf69daeadd4e4e4b8151ed888dfec20fb01728d89d56b3f38f2ae9c8c5, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413f, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd036413e},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{116, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h44ad339afbc21e9abf7b602a5ca535ea378135b6d10d81310bdd8293d1df3252, 264'h00b63ff7d0774770f8fe1d1722fa83acd02f434e4fc110a0cc8f6dddd37d56c463, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3e9a7582886089c62fb840cf3b83061cd1cff3ae4341808bb5bdee6191174177},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{117, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1260c2122c9e244e1af5151bede0c3ae23b54d7c596881d3eebad21f37dd878c, 256'h5c9a0c1a9ade76737a8811bd6a7f9287c978ee396aa89c11e47229d2ccb552f0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h24238e70b431b1a64efdf9032669939d4b77f249503fc6905feb7540dea3e6d2},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{118, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1877045be25d34a1d0600f9d5c00d0645a2a54379b6ceefad2e6bf5c2a3352ce, 264'h00821a532cc1751ee1d36d41c3d6ab4e9b143e44ec46d73478ea6a79a5c0e54159, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{119, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1877045be25d34a1d0600f9d5c00d0645a2a54379b6ceefad2e6bf5c2a3352ce, 264'h00821a532cc1751ee1d36d41c3d6ab4e9b143e44ec46d73478ea6a79a5c0e54159, 8'h01, 8'h01},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{120, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h455439fcc3d2deeceddeaece60e7bd17304f36ebb602adf5a22e0b8f1db46a50, 264'h00aec38fb2baf221e9a8d1887c7bf6222dd1834634e77263315af6d23609d04f77, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000002},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{121, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h455439fcc3d2deeceddeaece60e7bd17304f36ebb602adf5a22e0b8f1db46a50, 264'h00aec38fb2baf221e9a8d1887c7bf6222dd1834634e77263315af6d23609d04f77, 8'h01, 8'h02},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=8b(1B), s=8b(1B)
  '{122, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2e1f466b024c0c3ace2437de09127fed04b706f94b19a21bb1c2acf35cece718, 256'h0449ae3523d72534e964972cfd3b38af0bddd9619e5af223e4d1a40f34cf9f1d, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'h0000000000000000000000000000000000000000000000000000000000000003},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{123, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2e1f466b024c0c3ace2437de09127fed04b706f94b19a21bb1c2acf35cece718, 256'h0449ae3523d72534e964972cfd3b38af0bddd9619e5af223e4d1a40f34cf9f1d, 8'h01, 8'h03},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=8b(1B), s=8b(1B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2e1f466b024c0c3ace2437de09127fed04b706f94b19a21bb1c2acf35cece718, 256'h0449ae3523d72534e964972cfd3b38af0bddd9619e5af223e4d1a40f34cf9f1d, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364142, 256'h0000000000000000000000000000000000000000000000000000000000000003},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00dda95d7b0698de5d2d0b4f0034dbe35b50f978fcc518a84abf9c99efd96a2530, 256'h5adc08d6a63dbe831ab99cd9146e3c4c45492ad19521612542256d6af60e7888, 256'h0000000000000000000000000000000000000000000000000000000000000001, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd04917c8},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{126, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h02ef4d6d6cfd5a94f1d7784226e3e2a6c0a436c55839619f38fb4472b5f9ee77, 256'h7eb4acd4eebda5cd72875ffd2a2f26229c2dc6b46500919a432c86739f3ae866, 256'h0000000000000000000000000000000000000000000000000000000000000101, 256'hc58b162c58b162c58b162c58b162c58a1b242973853e16db75c8a1a71da4d39d},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{127, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h464f4ff715729cae5072ca3bd801d3195b67aec65e9b01aad20a2943dcbcb584, 264'h00b1afd29d31a39a11d570aa1597439b3b2d1971bf2f1abf15432d0207b10d1d08, 256'h000000000000000000000000000000000000000000000000002d9b4d347952cc, 256'hfcbc5103d0da267477d1791461cf2aa44bf9d43198f79507bd8779d69a13108e},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{128, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h157f8fddf373eb5f49cfcf10d8b853cf91cbcd7d665c3522ba7dd738ddb79a4c, 264'h00deadf1a5c448ea3c9f4191a8999abfcc757ac6d64567ef072c47fec613443b8f, 256'h000000000000000000000000000000000000001033e67e37b32b445580bf4efc, 256'h906f906f906f906f906f906f906f906ed8e426f7b1968c35a204236a579723d2},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{129, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h0934a537466c07430e2c48feb990bb19fb78cecc9cee424ea4d130291aa237f0, 264'h00d4f92d23b462804b5b68c52558c01c9996dbf727fccabbeedb9621a400535afa, 256'h0000000000000000000000000000000000000000000000000000000000000101, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{130, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d6ef20be66c893f741a9bf90d9b74675d1c2a31296397acb3ef174fd0b300c65, 256'h4a0c95478ca00399162d7f0f2dc89efdc2b28a30fbabe285857295a4b0c4e265, 256'h00000000000000000000000000000000000000062522bbd3ecbe7c39e93e7c26, 256'h783266e90f43dafe5cd9b3b0be86de22f9de83677d0f50713a468ec72fcf5d57},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{131, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00b7291d1404e0c0c07dab9372189f4bd58d2ceaa8d15ede544d9514545ba9ee06, 256'h29c9a63d5e308769cc30ec276a410e6464a27eeafd9e599db10f053a4fe4a829, 256'hfffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd03640c1, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{132, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00bb79f61857f743bfa1b6e7111ce4094377256969e4e15159123d9548acc3be6c, 256'h1f9d9f8860dcffd3eb36dd6c31ff2e7226c2009c4c94d8d7d2b5686bf7abd677, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h0000000000000000000000000000000000000000000000000000000000000001},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00bb79f61857f743bfa1b6e7111ce4094377256969e4e15159123d9548acc3be6c, 256'h1f9d9f8860dcffd3eb36dd6c31ff2e7226c2009c4c94d8d7d2b5686bf7abd677, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c1, 256'h0000000000000000000000000000000000000000000000000000000000000000},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{134, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d533b789a4af890fa7a82a1fae58c404f9a62a50b49adafab349c513b4150874, 256'h01b4171b803e76b34a9861e10f7bc289a066fd01bd29f84c987a10a5fb18c2d4, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{135, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3a3150798c8af69d1e6e981f3a45402ba1d732f4be8330c5164f49e10ec555b4, 256'h221bd842bc5e4d97eff37165f60e3998a424d72a450cf95ea477c78287d0343a, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{136, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3b37df5fb347c69a0f17d85c0c7ca83736883a825e13143d0fcfc8101e851e80, 256'h0de3c090b6ca21ba543517330c04b12f948c6badf14a63abffdf4ef8c7537026, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a0, 256'h7fffffffffffffffffffffffffffffff5d576e7357a4501ddfe92f46681b20a1},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{137, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00feb5163b0ece30ff3e03c7d55c4380fa2fa81ee2c0354942ff6f08c99d0cd82c, 264'h00e87de05ee1bda089d3e4e248fa0f721102acfffdf50e654be281433999df897e, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{138, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h238ced001cf22b8853e02edc89cbeca5050ba7e042a7a77f9382cd4149228976, 256'h40683d3094643840f295890aa4c18aa39b41d77dd0fb3bb2700e4f9ec284ffc2, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h44a5ad0bd0636d9e12bc9e0a6bdd5e1bba77f523842193b3b82e448e05d5f11e},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{139, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00961cf64817c06c0e51b3c2736c922fde18bd8c4906fcd7f5ef66c4678508f35e, 264'h00d2c5d18168cfbe70f2f123bd7419232bb92dd69113e2941061889481c5a027bf, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{140, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h13681eae168cd4ea7cf2e2a45d052742d10a9f64e796867dbdcb829fe0b10288, 256'h16528760d177376c09df79de39557c329cc1753517acffe8fa2ec298026b8384, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215b8, 256'haaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa9d1c9e899ca306ad27fe1945de0242b89},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{141, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5aa7abfdb6b4086d543325e5d79c6e95ce42f866d2bb84909633a04bb1aa31c2, 264'h0091c80088794905e1da33336d874e2f91ccf45cc59185bede5dd6f3f7acaae18b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'he91e1ba6ba898620a46bcb51dc0b8b4ad1dc35dad892c4552d1847b2ce444637},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{142, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 248'h277791b305a45b2b39590b2f05d3392a6c8182cef4eb540120e0f5c206c3e4, 256'h64108233fb0b8c3ac892d79ef8e0fbf92ed133addb4554270132584dc52eef41, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'he36bf0cec06d9b841da81332812f74f30bbaec9f202319206c6f0b8a0a400ff7},  // lens: hash=256b(32B), x=248b(31B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{143, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6efa092b68de9460f0bcc919005a5f6e80e19de98968be3cd2c770a9949bfb1a, 264'h00c75e6e5087d6550d5f9beb1e79e5029307bc255235e2d5dc99241ac3ab886c49, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'hea26b57af884b6c06e348efe139c1e4e9ec9518d60c340f6bac7d278ca08d8a6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{144, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h72d4a19c4f9d2cf5848ea40445b70d4696b5f02d632c0c654cc7d7eeb0c6d058, 264'h00e8c4cd9943e459174c7ac01fa742198e47e6c19a6bdb0c4f6c237831c1b3f942, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5b1d27a7694c146244a5ad0bd0636d9d9ef3b9fb58385418d9c982105077d1b7},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{145, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2a8ea2f50dcced0c217575bdfa7cd47d1c6f100041ec0e35512794c1be7e7402, 256'h58f8c17122ed303fda7143eb58bede70295b653266013b0b0ebd3f053137f6ec, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'hd27a7694c146244a5ad0bd0636d9e12abe687897e8e9998ddbd4e59a78520d0f},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{146, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0088de689ce9af1e94be6a2089c8a8b1253ffdbb6c8e9c86249ba220001a4ad3b8, 256'h0c4998e54842f413b9edb1825acbb6335e81e4d184b2b01c8bebdc85d1f28946, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'ha4f4ed29828c4894b5a17a0c6db3c256c2221449228a92dff7d76ca8206dd8dd},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{147, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00fea2d31f70f90d5fb3e00e186ac42ab3c1615cee714e0b4e1131b3d4d8225bf7, 264'h00b037a18df2ac15343f30f74067ddf29e817d5f77f8dce05714da59c094f0cda9, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h694c146244a5ad0bd0636d9e12bc9e09e60e68b90d0b5e6c5dddd0cb694d8799},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{148, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h7258911e3d423349166479dbe0b8341af7fbd03d0a7e10edccb36b6ceea5a3db, 256'h17ac2b8992791128fa3b96dc2fbd4ca3bfa782ef2832fc6656943db18e7346b0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h3d7f487c07bfc5f30846938a3dcef696444707cf9677254a92b06c63ab867d22},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{149, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h4f28461dea64474d6bb34d1499c97d37b9e95633df1ceeeaacd45016c98b3914, 264'h00c8818810b8cc06ddb40e8a1261c528faa589455d5a6df93b77bc5e0e493c7470, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6c7648fc0fbf8a06adb8b839f97b4ff7a800f11b1e37c593b261394599792ba4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{150, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h74f2a814fb5d8eca91a69b5e60712732b3937de32829be974ed7b68c5c2f5d66, 264'h00eff0f07c56f987a657f42196205f588c0f1d96fd8a63a5f238b48f478788fe3b, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h9be363a286f23f6322c205449d320baad417953ecb70f6214e90d49d7d1f26a8},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{151, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h195b51a7cc4a21b8274a70a90de779814c3c8ca358328208c09a29f336b82d6a, 264'h00b2416b7c92fffdc29c3b1282dd2a77a4d04df7f7452047393d849989c5cee9ad, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h29798c5c45bdf58b4a7b2fdc2c46ab4af1218c7eeb9f0f27a88f1267674de3b0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{152, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h622fc74732034bec2ddf3bc16d34b3d1f7a327dd2a8c19bab4bb4fe3a24b58aa, 256'h736b2f2fae76f4dfaecc9096333b01328d51eb3fda9c9227e90d0b449983c4f0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h0b70f22ca2bb3cefadca1a5711fa3a59f4695385eb5aedf3495d0b6d00f8fd85},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{153, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1f7f85caf2d7550e7af9b65023ebb4dce3450311692309db269969b834b611c7, 256'h0827f45b78020ecbbaf484fdd5bfaae6870f1184c21581baf6ef82bd7b530f93, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h16e1e459457679df5b9434ae23f474b3e8d2a70bd6b5dbe692ba16da01f1fb0a},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{154, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h49c197dc80ad1da47a4342b93893e8e1fb0bb94fc33a83e783c00b24c781377a, 264'h00efc20da92bac762951f72474becc734d4cc22ba81b895e282fdac4df7af0f37d, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2252d685e831b6cf095e4f0535eeaf0ddd3bfa91c210c9d9dc17224702eaf88f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{155, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00d8cb68517b616a56400aa3868635e54b6f699598a2f6167757654980baf6acbe, 256'h7ec8cf449c849aa03461a30efada41453c57c6e6fbc93bbc6fa49ada6dc0555c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h75135abd7c425b60371a477f09ce0f274f64a8c6b061a07b5d63e93c65046c53},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{156, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h030713fb63f2aa6fe2cadf1b20efc259c77445dafa87dac398b84065ca347df3, 264'h00b227818de1a39b589cb071d83e5317cccdc2338e51e312fe31d8dc34a4801750, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'hd55555555555555555555555555555547c74934474db157d2a8c3f088aced62a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{157, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00babb3677b0955802d8e929a41355640eaf1ea1353f8a771331c4946e3480afa7, 256'h252f196c87ed3d2a59d3b1b559137fed0013fecefc19fb5a92682b9bca51b950, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'hc1777c8853938e536213c02464a936000ba1e21c0fc62075d46c624e23b52f31},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{158, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1aab2018793471111a8a0e9b143fde02fc95920796d3a63de329b424396fba60, 264'h00bbe4130705174792441b318d3aa31dfe8577821e9b446ec573d272e036c4ebe9, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h30bbb794db588363b40679f6c182a50d3ce9679acdd3ffbe36d7813dacbdc818},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{159, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008cb0b909499c83ea806cd885b1dd467a0119f06a88a0276eb0cfda274535a8ff, 256'h47b5428833bc3f2c8bf9d9041158cf33718a69961cd01729bc0011d1e586ab75, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2c37fd995622c4fb7fffffffffffffffc7cee745110cb45ab558ed7c90c15a2f},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{160, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008f03cf1a42272bb1532723093f72e6feeac85e1700e9fbe9a6a2dd642d74bf5d, 256'h3b89a7189dad8cf75fc22f6f158aa27f9c2ca00daca785be3358f2bda3862ca0, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h7fd995622c4fb7ffffffffffffffffff5d883ffab5b32652ccdcaa290fccb97d},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{161, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h44de3b9c7a57a8c9e820952753421e7d987bb3d79f71f013805c897e018f8ace, 264'h00a2460758c8f98d3fdce121a943659e372c326fff2e5fc2ae7fa3f79daae13c12, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'hffb32ac4589f6ffffffffffffffffffebb107ff56b664ca599b954521f9972fa},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{162, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h6fb8b2b48e33031268ad6a517484dc8839ea90f6669ea0c7ac3233e2ac31394a, 256'h0ac8bbe7f73c2ff4df9978727ac1dfc2fd58647d20f31f99105316b64671f204, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h5622c4fb7fffffffffffffffffffffff928a8f1c7ac7bec1808b9f61c01ec327},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{163, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00bea71122a048693e905ff602b3cf9dd18af69b9fc9d8431d2b1dd26b942c95e6, 264'h00f43c7b8b95eb62082c12db9dbda7fe38e45cbe4a4886907fb81bdb0c5ea9246c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h44104104104104104104104104104103b87853fd3b7d3f8e175125b4382f25ed},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{164, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00da918c731ba06a20cb94ef33b778e981a404a305f1941fe33666b45b03353156, 264'h00e2bb2694f575b45183be78e5c9b5210bf3bf488fd4c8294516d89572ca4f5391, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2739ce739ce739ce739ce739ce739ce705560298d1f2f08dc419ac273a5b54d9},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{165, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3007e92c3937dade7964dfa35b0eff031f7eb02aed0a0314411106cdeb70fe3d, 256'h5a7546fc0552997b20e3d6f413e75e2cb66e116322697114b79bac734bfc4dc5, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'hb777777777777777777777777777777688e6a1fe808a97a348671222ff16b863},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{166, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h60e734ef5624d3cbf0ddd375011bd663d6d6aebc644eb599fdf98dbdcd18ce9b, 264'h00d2d90b3ac31f139af832cccf6ccbbb2c6ea11fa97370dc9906da474d7d8a7567, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h6492492492492492492492492492492406dd3a19b8d5fb875235963c593bd2d3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{167, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0085a900e97858f693c0b7dfa261e380dad6ea046d1f65ddeeedd5f7d8af0ba337, 256'h69744d15add4f6c0bc3b0da2aec93b34cb8c65f9340ddf74e7b0009eeeccce3c, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h955555555555555555555555555555547c74934474db157d2a8c3f088aced62c},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{168, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h38066f75d88efc4c93de36f49e037b234cc18b1de5608750a62cab0345401046, 264'h00a3e84bed8cfcb819ef4d550444f2ce4b651766b69e2e2901f88836ff90034fed, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h2aaaaaaaaaaaaaaaaaaaaaaaaaaaaaaa3e3a49a23a6d8abe95461f8445676b17},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{169, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h0098f68177dc95c1b4cbfa5245488ca523a7d5629470d035d621a443c72f39aabf, 264'h00a33d29546fa1c648f2c7d5ccf70cf1ce4ab79b5db1ac059dbecd068dbdff1b89, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'hbffffffffffffffffffffffffffffffebaaedce6af48a03bbfd25e8cd0364143},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{170, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h5c2bbfa23c9b9ad07f038aa89b4930bf267d9401e4255de9e8da0a5078ec8277, 264'h00e3e882a31d5e6a379e0793983ccded39b95c4353ab2ff01ea5369ba47b0c3191, 256'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffc, 256'h185ddbca6dac41b1da033cfb60c152869e74b3cd66e9ffdf1b6bc09ed65ee40c},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{171, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2ea7133432339c69d27f9b267281bd2ddd5f19d6338d400a05cd3647b157a385, 256'h3547808298448edb5e701ade84cd5fb1ac9567ba5e8fb68a6b933ec4b5cc84cc, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 256'hd612c2984c2afa416aa7f2882a486d4a8426cb6cfc91ed5b737278f9fca8be68},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2ea7133432339c69d27f9b267281bd2ddd5f19d6338d400a05cd3647b157a385, 264'h00cab87f7d67bb7124a18fe5217b32a04e536a9845a1704975946cc13a4a337763, 256'h32b0d10d8d0e04bc8d4d064d270699e87cffc9b49c5c20730e1c26f6105ddcda, 256'hd612c2984c2afa416aa7f2882a486d4a8426cb6cfc91ed5b737278f9fca8be68},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{173, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008aa2c64fa9c6437563abfbcbd00b2048d48c18c152a2a6f49036de7647ebe82e, 256'h1ce64387995c68a060fa3bc0399b05cc06eec7d598f75041a4917e692b7f51ff, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0, 256'h33333333333333333333333333333332f222f8faefdb533f265d461c29a47373},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{174, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h391427ff7ee78013c14aec7d96a8a062209298a783835e94fd6549d502fff71f, 264'h00dd6624ec343ad9fcf4d9872181e59f842f9ba4cccae09a6c0972fb6ac6b4c6bd, 256'hc6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{175, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00e762b8a219b4f180219cc7a9059245e4961bd191c03899789c7a34b89e8c138e, 264'h00c1533ef0419bb7376e0bfde9319d10a06968791d9ea0eed9c1ce6345aed9759e, 256'hc6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'hb6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{176, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h009aedb0d281db164e130000c5697fae0f305ef848be6fffb43ac593fbb950e952, 264'h00fa6f633359bdcd82b56b0b9f965b037789d46b9a8141b791b2aefa713f96c175, 256'hc6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h99999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{177, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008ad445db62816260e4e687fd1884e48b9fc0636d031547d63315e792e19bfaee, 256'h1de64f99d5f1cd8b6ec9cb0f787a654ae86993ba3db1008ef43cff0684cb22bd, 256'hc6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{178, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h1f5799c95be89063b24f26e40cb928c1a868a76fb0094607e8043db409c91c32, 264'h00e75724e813a4191e3a839007f08e2e897388b06d4a00de6de60e536d91fab566, 256'hc6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{179, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00a3331a4e1b4223ec2c027edd482c928a14ed358d93f1d4217d39abf69fcb5ccc, 256'h28d684d2aaabcd6383775caa6239de26d4c6937bb603ecb4196082f4cffd509d, 256'hc6047f9441ed7d6d3045406e95c07cd85c778e4b8cef3ca7abac09b95c709ee5, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{180, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h3f3952199774c7cf39b38b66cb1042a6260d8680803845e4d433adba3bb24818, 256'h5ea495b68cbc7ed4173ee63c9042dc502625c7eb7e21fb02ca9a9114e0a3a18d, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h55555555555555555555555555555554e8e4f44ce51835693ff0ca2ef01215c0},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{181, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00cdfb8c0f422e144e137c2412c86c171f5fe3fa3f5bbb544e9076288f3ced786e, 256'h054fd0721b77c11c79beacb3c94211b0a19bda08652efeaf92513a3b0a163698, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'hb6db6db6db6db6db6db6db6db6db6db5f30f30127d33e02aad96438927022e9c},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{182, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h73598a6a1c68278fa6bfd0ce4064e68235bc1c0f6b20a928108be336730f87e3, 264'h00cbae612519b5032ecc85aed811271a95fe7939d5d3460140ba318f4d14aba31d, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h99999999999999999999999999999998d668eaf0cf91f9bd7317d2547ced5a5a},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{183, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h58debd9a7ee2c9d59132478a5440ae4d5d7ed437308369f92ea86c82183f10a1, 256'h6773e76f5edbf4da0e4f1bdffac0f57257e1dfa465842931309a24245fda6a5d, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h66666666666666666666666666666665e445f1f5dfb6a67e4cba8c385348e6e7},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{184, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h008b904de47967340c5f8c3572a720924ef7578637feab1949acb241a5a6ac3f5b, 264'h00950904496f9824b1d63f3313bae21b89fae89afdfc811b5ece03fd5aa301864f, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h49249249249249249249249249249248c79facd43214c011123c1b03a93412a5},  // lens: hash=256b(32B), x=264b(33B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{185, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 264'h00f4892b6d525c771e035f2a252708f3784e48238604b4f94dc56eaa1e546d941a, 256'h346b1aa0bce68b1c50e5b52f509fb5522e5c25e028bc8f863402edb7bcad8b1b, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h0eb10e5ab95f2f275348d82ad2e4d7949c8193800d8c9c75df58e343f0ebba7b},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{186, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{187, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 256'h483ada7726a3c4655da4fbfc0e1108a8fd17b448a68554199c47d08ffb10d4b8, 256'h44a5ad0bd0636d9e12bc9e0a6bdd5e1bba77f523842193b3b82e448e05d5f11e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{188, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{189, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h79be667ef9dcbbac55a06295ce870b07029bfcdb2dce28d959f2815b16f81798, 264'h00b7c52588d95c3b9aa25b0403f1eef75702e84bb7597aabe663b82f6f04ef2777, 256'h44a5ad0bd0636d9e12bc9e0a6bdd5e1bba77f523842193b3b82e448e05d5f11e, 256'h2492492492492492492492492492492463cfd66a190a6008891e0d81d49a0952},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{190, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'hf80ae4f96cdbc9d853f83d47aae225bf407d51c56b7776cd67d0dc195d99a9dc, 256'hb303e26be1f73465315221f0b331528807a1a9b6eb068ede6eebeaaa49af8a36},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{191, 1'b1, 256'hdc1921946f4af96a2856e7be399007c9e807bdf4c5332f19f59ec9dd1bb8c7b3, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h109cd8ae0374358984a8249c0a843628f2835ffad1df1a9a69aa2fe72355545c, 256'hac6f00daf53bd8b1e34da329359b6e08019c5b037fed79ee383ae39f85a159c6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{192, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'hd035ee1f17fdb0b2681b163e33c359932659990af77dca632012b30b27a057b3, 256'h1939d9f3b2858bc13e3474cb50e6a82be44faa71940f876c1cba4c3e989202b6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{193, 1'b1, 256'hde47c9b27eb8d300dbb5f2c353e632c393262cf06340c4fa7f1b40c4cbd36f90, 256'h782c8ed17e3b2a783b5464f33b09652a71c678e05ec51e84e2bcfc663a3de963, 264'h00af9acb4280b8c7f7c42f4ef9aba6245ec1ec1712fd38a0fa96418d8cd6aa6152, 256'h4f053f563ad34b74fd8c9934ce59e79c2eb8e6eca0fef5b323ca67d5ac7ed238, 256'h4d4b05daa0719e773d8617dce5631c5fd6f59c9bdc748e4b55c970040af01be5},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{194, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h6d6a4f556ccce154e7fb9f19e76c3deca13d59cc2aeb4ecad968aab2ded45965, 256'h53b9fa74803ede0fc4441bf683d56c564d3e274e09ccf47390badd1471c05fb7},  // lens: hash=256b(32B), x=256b(32B), y=232b(29B), r=256b(32B), s=256b(32B)
  '{195, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'haad503de9b9fd66b948e9acf596f0a0e65e700b28b26ec56e6e45e846489b3c4, 256'hfff223c5d0765447e8447a3f9d31fd0696e89d244422022ff61a110b2a8c2f04},  // lens: hash=256b(32B), x=256b(32B), y=232b(29B), r=256b(32B), s=256b(32B)
  '{196, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 232'h01060492d5a5673e0f25d8d50fb7e58c49d86d46d4216955e0aa3d40e1, 256'h9182cebd3bb8ab572e167174397209ef4b1d439af3b200cdf003620089e43225, 256'habb88367d15fe62d1efffb6803da03109ee22e90bc9c78e8b4ed23630b82ea9d},  // lens: hash=256b(32B), x=256b(32B), y=232b(29B), r=256b(32B), s=256b(32B)
  '{197, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h3854a3998aebdf2dbc28adac4181462ccac7873907ab7f212c42db0e69b56ed8, 256'hc12c09475c772fd0c1b2060d5163e42bf71d727e4ae7c03eeba954bf50b43bb3},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{198, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'he94dbdc38795fe5c904d8f16d969d3b587f0a25d2de90b6d8c5c53ff887e3607, 256'h856b8c963e9b68dade44750bf97ec4d11b1a0a3804f4cb79aa27bdea78ac14e4},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{199, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6e823555452914099182c6b2c1d6f0b5d28d50ccd005af2ce1bba541aa40caff, 264'h00fffffffef9fb6d2a5a98c1f0da272af0481a73b62792b92bde96aa1e55c2bb4e, 256'h49fc102a08ca47b60e0858cd0284d22cddd7233f94aaffbb2db1dd2cf08425e1, 256'h5b16fca5a12cdb39701697ad8e39ffd6bdec0024298afaa2326aea09200b14d6},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{200, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h41efa7d3f05a0010675fcb918a45c693da4b348df21a59d6f9cd73e0d831d67a, 256'hbbab52596c1a1d9484296cdc92cbf07e665259a13791a8fe8845e2c07cf3fc67},  // lens: hash=256b(32B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{201, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'hb615698c358b35920dd883eca625a6c5f7563970cdfc378f8fe0cee17092144c, 256'hda0b84cd94a41e049ef477aeac157b2a9bfa6b7ac8de06ed3858c5eede6ddd6d},  // lens: hash=256b(32B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{202, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h013fd22248d64d95f73c29b48ab48631850be503fd00f8468b5f0f70e0, 264'h00f6ee7aa43bc2c6fd25b1d8269241cbdd9dbb0dac96dc96231f430705f838717d, 256'h87cf8c0eb82d44f69c60a2ff5457d3aaa322e7ec61ae5aecfd678ae1c1932b0e, 256'hc522c4eea7eafb82914cbf5c1ff76760109f55ddddcf58274d41c9bc4311e06e},  // lens: hash=256b(32B), x=232b(29B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{203, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'h62f48ef71ace27bf5a01834de1f7e3f948b9dce1ca1e911d5e13d3b104471d82, 256'ha1570cc0f388768d3ba7df7f212564caa256ff825df997f21f72f5280d53011f},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{204, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'hf6b0e2f6fe020cf7c0c20137434344ed7add6c4be51861e2d14cbda472a6ffb4, 256'h9be93722c1a3ad7d4cf91723700cb5486de5479d8c1b38ae4e8e5ba1638e9732},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{205, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h25afd689acabaed67c1f296de59406f8c550f57146a0b4ec2c97876dffffffff, 264'h00fa46a76e520322dfbc491ec4f0cc197420fc4ea5883d8f6dd53c354bc4f67c35, 256'hdb09d8460f05eff23bc7e436b67da563fa4b4edb58ac24ce201fa8a358125057, 256'h46da116754602940c8999c8d665f786c50f5772c0a3cdbda075e77eabc64df16},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{206, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'h592c41e16517f12fcabd98267674f974b588e9f35d35406c1a7bb2ed1d19b7b8, 256'hc19a5f942607c3551484ff0dc97281f0cdc82bc48e2205a0645c0cf3d7f59da0},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{207, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'hbe0d70887d5e40821a61b68047de4ea03debfdf51cdf4d4b195558b959a032b2, 256'h8266b4d270e24414ecacb14c091a233134b918d37320c6557d60ad0a63544ac4},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{208, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 264'h00d12e6c66b67734c3c84d2601cf5d35dc097e27637f0aca4a4fdb74b6aadd3bb9, 256'h3f5bdff88bd5736df898e699006ed750f11cf07c5866cd7ad70c7121ffffffff, 256'hfae92dfcb2ee392d270af3a5739faa26d4f97bfd39ed3cbee4d29e26af3b206a, 256'h93645c80605595e02c09a0dc4b17ac2a51846a728b3e8d60442ed6449fd3342b},  // lens: hash=256b(32B), x=264b(33B), y=256b(32B), r=256b(32B), s=256b(32B)
  '{209, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h176a2557566ffa518b11226694eb9802ed2098bfe278e5570fe1d5d7af18a943, 256'hed6e2095f12a03f2eaf6718f430ec5fe2829fd1646ab648701656fd31221b97d},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{210, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'h60be20c3dbc162dd34d26780621c104bbe5dace630171b2daef0d826409ee5c2, 256'hbd8081b27762ab6e8f425956bf604e332fa066a99b59f87e27dc1198b26f5caa},  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
  '{211, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 256'h6d4a7f60d4774a4f0aa8bbdedb953c7eea7909407e3164755664bc2800000000, 264'h00e659d34e4df38d9e8c9eaadfba36612c769195be86c77aac3f36e78b538680fb, 256'hedf03cf63f658883289a1a593d1007895b9f236d27c9c1f1313089aaed6b16ae, 256'he5b22903f7eb23adc2e01057e39b0408d495f694c83f306f1216c9bf87506074}  // lens: hash=256b(32B), x=256b(32B), y=264b(33B), r=256b(32B), s=256b(32B)
};
`endif // WYCHERPROOF_SECP256K1_SHA256_P1363_SV
