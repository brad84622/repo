`ifndef WYCHERPROOF_SECP224R1_SHA256_SV
`define WYCHERPROOF_SECP224R1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp224r1_sha256;

localparam int TEST_VECTORS_SECP224R1_SHA256_NUM = 73;

ecdsa_vector_secp224r1_sha256 test_vectors_secp224r1_sha256 [] = '{
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{113, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 0, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=0b(0B), s=224b(28B)
  '{114, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 0},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=0b(0B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h38de5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{118, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h637d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{119, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a84, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{120, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad901},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{121, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=216b(27B), s=224b(28B)
  '{122, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 216'hde5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=216b(27B), s=224b(28B)
  '{123, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 216'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad9},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=216b(27B)
  '{124, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 216'h7d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=216b(27B)
  '{129, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=224b(28B)
  '{130, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=8b(1B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'hc521a3f9db5a98812849baf26bdf441fd72b663dc4161062747575fc, 224'h617d6af141efd0c800c9ba3382c2faf758540a5dd98d1756a1dad981},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{140, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h3ade5c0624a5677ed7b6450d9420bbe028d499c23be9ef9d8b8a8a04, 224'h9e82950ebe102f37ff3645cc7d3d0508a7abf5a22672e8a95e25267f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{144, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{145, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{146, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h00, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{154, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{155, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{156, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'h01, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{164, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{165, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{166, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 8'hff, 8'hff},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{232, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h59a9f83289ef6995d5d5592e80ab4f6a81123f69d385d3cfb152faf2, 224'h3a97d5be190d5819241067e2be56375ab84155baab8fc7aeb7f8cb3d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{241, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h5984af8c89fb9d596a1f28fd3d41e46f7205fe12fa63437ac79e7e81, 224'h33b16b742d45f18f88de2713078384e6150f06b8b99f36ab2ce3dd49},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{248, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4769fba554fd436051c285bdadfa33a443d4f7084dd598ce3b98b8fb, 224'h0c014c87cb14113d75864f74905f75b34f9970ba58b5d0676021826d},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{258, 1'b1, 256'h3760a7f37cf96218f29ae43732e513efd2b6f552ea4b6895464b9300000000c8, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h0a1c2c2478e244464226c660edf724db1213f4923eb725d611d976fd, 224'h764e55186a76f734891d05fb57af2727fab8fbea684ca4321d5de540},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{269, 1'b1, 256'hde030419345ca15c75ffffffff8074799b9e0956cc43135d16dfbe4d27d7e68d, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h1b393477941879271873a8c043a77caadb9957fcdd263a6ac978e4ba, 224'h270060d5f356ebb6d185772baa78b878af6807378e0d5c532da0a4a7},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{273, 1'b1, 256'hac18f8418c55a2502cb7d53f9affffffff5c31d89fda6a6b8476397c04edf411, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h74a4c51dd60c7118467be29652060f39af94f8c0eb7f15c64771010c, 224'h6102ec0c9257e607af3f3ff7490b54e78111f422bec11ba01277171f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{281, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h7e0f48761089aa4c7ecd5a7ac5380836b1e5d381d3400174d15df98b, 224'h0c3df50060e3a6714aa565a33d784e7b16ac87bebfb3c2255cfd832c},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{282, 1'b1, 256'h1273b4502ea4e3bccee044ee8e8db7f774ecbcd52e8ceb571757ffffffffe20a, 232'h00eada93be10b2449e1e8bb58305d52008013c57107c1a20a317a6cba7, 232'h00eca672340c03d1d2e09663286691df55069fa25490c9dd9f9c0bb2b5, 224'h4d6f7408508eb0814dcd48007f0efd9e2b91cdac4030540cc678de19, 224'h1e74f8dc34d13613ef42462fe88981cbe2489be10e4cdae975a1b38e},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{289, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h20888e1c0f5694c4c0363b36482beb6e1e6649b3d3b26f127febb6fc, 232'h00de00c2f3d8e4a7e8a0bafd417c96d3e81c975946a2f3686aa39d35f1, 224'h7fffffffffffffffffffffffffffffffffffffffffffffffffffffff, 224'h3d5052691b8dc89debad360466f2a39e82e8ae2aefb77c3c92ad7cd1},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{291, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h579d53f39d5109bd440e3e3e7efd603740963348ff9c72c03b0fe6b8, 232'h00df02f133ecd60b072a0812adc752708f2be9d8c9ad5953d8c7bf3965, 8'h03, 8'h01},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{292, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d2a14c8106d89f3536faebdafcd4680f65ab4bf2243164ca1464b628, 232'h00acaf2bee52e6231d3c980f52f8e189a41c3e3a05e591195ec864217a, 8'h03, 8'h03},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=8b(1B), s=8b(1B)
  '{293, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00e892479153ad13ea5ca45d4c323ebf1fc3cd0cdf787c34306a3f79a4, 224'h326ca9645f2b517608dc1f08b7a84cfc61e6ff68d14f27d2043c7ef5, 8'h03, 8'h04},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=8b(1B), s=8b(1B)
  '{297, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00f293a8a2b4aff0bed95c663b364afe69778d38dd7e7a304f7d3c74e6, 224'h17dfd09e7803c4439a6c075cb579cde652d03f7559ff58846312fa4c, 56'h2d9b4d347952cc, 224'h3e85d56474b5c55fbe86608442a84b2bf093b7d75f53a47250e1c70c},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=56b(7B), s=224b(28B)
  '{298, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d4ddf003b298cbaa7d2edc584b28b474a76162ed4b5b0f6222c54317, 232'h00d4e4fe030f178fb4aa4a6d7f61265ecd7ef13c313606b8d341a8b954, 104'h1033e67e37b32b445580bf4efb, 224'h02fd02fd02fd02fd02fd02fd02fd0043a4fd2da317247308c74dc6b8},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=104b(13B), s=224b(28B)
  '{302, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a7f7b99e5cdc6fec8928eff773ccdf3b68b19d43cdb41809e19c60f3, 224'h1736b7a0c12a9c2d706671912915142b3e05c89ef3ad497bd6c34699, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h01},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{303, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a7f7b99e5cdc6fec8928eff773ccdf3b68b19d43cdb41809e19c60f3, 224'h1736b7a0c12a9c2d706671912915142b3e05c89ef3ad497bd6c34699, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 8'h00},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=8b(1B)
  '{304, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h009cf00010b4ad86636f6cc70fb58c3b995c0d12e46fc58e24b0d28f69, 224'h21c8a8a320cc450ccb15ebd71617f4ed25db4d3413fbdf157d31dbb6, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00ae9b3636b8547232df438559b5a109e0238a73a76afc25d070ea2742, 224'h7210a69de44ad645b1b03845040f46fce238e92c131a71e4b184c01f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008d57d4fce62757791888c1938076fd766daeb2ec9f1bda8ad5df4809, 232'h00aade924d7ea3ae5abbd0719a7d4865759da654cf76cf7ec031277108, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f, 224'h7fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e151f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{308, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h008a5dfedc9dd1cb9a439c88b3dd472b2e66173f7866855db6bb6c12fd, 224'h3badfbb8a4c6fd80e66510957927c78a2aa02ecef62816d0356b49c3, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h44a5ad0bd0636d9e12bc9e0a6bdc74bfe082087ae8b61cbd54b8103f},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{309, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h0083a59fc3df295e84c290b32d0b550a06f99456fc2298e4a68c4f2bff, 224'h1b34f483db30db3a51d8288732c107d8b1a858cd54c3936e1b5c11a4, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{314, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h44e309eb686e7af7f1e2cc17fd56542b38910b3b7908ea54fb038d36, 224'h477e829d4c8332e5b29f344ad27a21c18dab24a31ce7985b63a21304, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h074aae944ee7a7d544a5ad0bd06366f872d2250ba3018a63d2a7f2e6},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{316, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00c46c1ad3d3d0df8e9c0f525c21ce8d81ef9d66297f442d6309966722, 224'h0cfa2253aa31a98d8966b85969bf9c819c019292ef6a53ac1db2a108, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h55d289dcf4faa894b5a17a0c6db3741bbc4ecbe01d01ea33ee7a4e7b},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b7b2e48c1e60e20925f4d9b6be600dd83786a936c9bfab00639c33ca, 232'h00a967cbc65070739a3379da80d54843a18d9c11a29a32234a0b303c12, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h4ee7a7d544a5ad0bd0636d9e12bc561ce04faaf1312bba3a15601ebc},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{318, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00f4a3d4598875af7f2741bbd67b1733b6541bc5325b3bcb4d3267c27e, 232'h00c30bf322f58a45c6c2aa2ced55f175d1cbf72a7c5bfc464d74f666c0, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h361b9cd74d65e79a5874c501bca4973b20347ec97f6de10072d8b46a},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h56d1e5c1d664f6ce2fc1fcb937a7ce231a29486abf36c73f77a2bd11, 224'h6cb282c9d7c6fc05f399c183e880ea362edf043cd28ffac9f94f2141, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c3739ae9acbcf34b0e98a0379492e764068fd92fedbc200e5b168d4},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{322, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h113a2cc57c8ee7de11bc45e14546c72a29725b9a7218114ac31f0281, 224'h6c765b9a46b0215312a3292f5979c98d37b35883baa156281b1bae8c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffffb2364ae85014b149b86c741eb8be},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00bbce4b17d45d24a1c80bc8eca98c359d5e1e458058a00b950643256d, 232'h00fe09e092318e39303dca03688e4ecf300300784312d617e5088c584c, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h2db5f61aea817276af2064e104c7a30e32034cb526dd0aacfa56566f},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00911c0033eac46332691cb7920c4950eed57354761e1081a1ea9f1279, 224'h508ebf7cfd3eab5dabdee1be14ce8296b1fc20acfaac16f7824c6002, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h6c7513e5f48c07ffffffffffffff9d21fd1b31544cb13ca86a75b25e},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{328, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h0f759330e7992752aae6a85f7bb0599784bea53e288ff7ee8d53d5e6, 232'h00defe617362380e92f9a23c4fdcc34e09713aab9cc44119418f6f2fd1, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3e5f48c07fffffffffffffffffffc724968c0ecf9ed783744a7337b3},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h2bcf4371b319a691ed0e2e0c4a55a8a9b987dec86b863621e97b9c09, 224'h5b8660a74cc964a6af0311edc6b1cd980f9c7bf3a6c9b7f9132a0b2f, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h7fffffffffffffffffffffffffff646c95d0a029629370d8e83d717f},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00a6f252568f6fbd1ae045e602344359c0c216911723748f9a3e7fadec, 224'h3b76efc75ba030bfe7de2ded686991e6183d40241a05b479693c7015, 224'h7ffffffffffffffffffffffffffffffffffffffffffffffffffffffd, 224'h3fffffffffffffffffffffffffff8b51705c781f09ee94a2ae2e1520},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{335, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h3672ba9718e60d00eab4295c819ea366a778dd6fd621fa9665259cb6, 224'h7ae5e847eeaea674beeb636379e968f79265502e414a1d444f04ae79, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h33eeefbfc77229136e56b575144863ed90b4c0f8a9e315816d6de648, 224'h051749dd11480c141fb5a1946313163c0141265b68a26216bcb9936a, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h5555555555555555555555555555078ba03da56a069f0dc1c9740e14},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{338, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h7abba0cbff134ddcf54d04846f954b882ca9faefdfe818898bfb378b, 224'h792f10b57970ae57bb4fb01c08886848855aeb1984d3d6fcb2b412df, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h33333333333333333333333333330486f9be9672d0c5d50ddf45a20c},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{340, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 224'h065d9ef133ce81c2d6b66e928360f9527f8f36b5badd35b5f1093427, 224'h2004852755f77440a0b08b9f165489c0696e8b4981d6d04a285b0fd1, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89852},  // lens: hash=256b(32B), x=224b(28B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{341, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00d6cea09472ede574ce1e0546c9acd0e1cd8cba9b121df29e89d5092e, 232'h0083904ebfb902ea61c987dc0508e0c9a7e563e2609feaf79140ab91d6, 224'h706a46dc76dcb76798e60e6d89474788d16dc18032d268fd1a704fa6, 224'h0eb10e5ab95facded4061029d63a46f46f12947411f2ea561a592057},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{349, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 232'h00bd376388b5f723fb4c22dfe6cd4375a05a07476444d5819985007e34, 224'h44a5ad0bd0636d9e12bc9e0a6bdc74bfe082087ae8b61cbd54b8103f, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{351, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 232'h00b70e0cbd6bb4bf7f321390b94a03c1d356c21122343280d6115c1d21, 224'h42c89c774a08dc04b3dd201932bc8a5ea5f8b89bbb2a7e667aff81cd, 224'h44a5ad0bd0636d9e12bc9e0a6bdc74bfe082087ae8b61cbd54b8103f, 224'h249249249249249249249249249227ce201a6b76951f982e7ae89851},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{356, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00aed6fcad2400c4d94e55dbb6b012ce3d4c2b46843fbe99d4289e6ecf, 232'h008a24a89e71343d7d151d258d2cb690349c2d56b366dd10a600000000, 224'h519bf185ff4635271961fa491be257231deeea9c53a6ede3b4a89ed1, 224'h486bdad484a6a3134e1471cf56a9df0fac50f773b3e37d6f327617d7},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{360, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h76be0112674ec29128823e1af7512e6143872fef30a64e2f1799bd56, 224'h187e503e1a48c27b549fe0a4ce5e581e242c8663fc9efb02d6f2b193},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{361, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00bf19ecfe43ffe289f699f479316145b9a7f7370b9ece5ab1212174f1, 224'h73d528949ae9142f818bade71a960407963be0b6482a6a60ffffffff, 224'h36245ef126b5b51e459f84eaaad5a495061f0471dc8c23f1c5f16282, 224'h39e31d72a06ba8e14fcf95778e07bc16a2628e39449da8857d506edc},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{362, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h26e5abf135cb54eaaa16b69e4b0b292275344e88a09df6df80000000, 232'h00eab891de54e3f26ff50ab989f333dac551583d468ae623c596434af0, 224'h258682975df8bca7f203f771ebeb478ef637360c860fc386cfb21745, 224'h7663e70188047e41469a2a35c8c330dd900f2340ba82aafd22962a96},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{365, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ec627f345545d03f8c6dbd08e575527116567fe375f9ecaaffffffff, 224'h41bf705697d5f716bcf78718d5393b63a98691f4a1f24246375538fd, 224'h19397fe5d3ecabf80fc624c1bf379564387517c185087dc97d605069, 224'h33b5773e9aaf6c34cb612cfc81efd3bf9c22224e8c4fa1bfccf5c501},  // lens: hash=256b(32B), x=232b(29B), y=224b(28B), r=224b(28B), s=224b(28B)
  '{372, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 224'h15016e52b36472d536477605fb805dd3903082a062d1ea30af9e555a, 232'h00ffffffff89d2d70e023de6e7b07e97df400a992b9a4a0e0ce178d20c, 224'h32fa0ca7e07f1f86ac350734994e1f31b6da9c82f93dced2b983c29c, 224'h7b7891282206a45711bdfcb2a102b5d289df84ff5778548603574004},  // lens: hash=256b(32B), x=224b(28B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{378, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h1f81cd924362ec825890307b9b3936e0d8f728a7c84bdb43c5cf0433, 224'h39d3e46a03040ad41ac026b18e0629f6145e3dc8d1e6bbe200c8482b},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{379, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00ffffffffeadf7cee8d34d04cf22c8f7de35674fb2f501d242a76f725, 232'h0086c409309d398e60ce1e0a4c9e05a9d32627577e8ce2cc7f3afa2c3e, 224'h00fda613aa67ca42673ad4309f3f0f05b2569f3dee63f4aa9cc54cf3, 224'h1e5a64b68a37e5b201c918303dc7a40439aaeacf019c5892a8f6d0ce},  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
  '{382, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 192'h0e2ab0e8495e859eb2afb00769d6e7fe626a119167c0b6bc, 224'h6e54f941204d4639b863c98a65b7bee318d51ab1900a8f345eac6f07, 224'h0da5054829214ecde5e10579b36a2fe6426c24b064ed77c38590f25c},  // lens: hash=256b(32B), x=232b(29B), y=192b(24B), r=224b(28B), s=224b(28B)
  '{385, 1'b1, 256'h2f77668a9dfbf8d5848b9eeb4a7145ca94c6ed9236e4a773f6dcafa5132b2f91, 232'h00b0013c6fbff6f09fecda1c263ef65399d4cf989ca5fc4f8fff0fe9e1, 232'h00fffffffff1d54f17b6a17a614d504ff7962918019d95ee6e983f4945, 224'h1526eb2f657ebea9af4ca184b975c02372c88e24e835f3f5774c0e12, 224'h1f1ecce38ee52372cb201907794de17b6d6c1afa13c316c51cb07bc7}  // lens: hash=256b(32B), x=232b(29B), y=232b(29B), r=224b(28B), s=224b(28B)
};
`endif // WYCHERPROOF_SECP224R1_SHA256_SV
