`ifndef WYCHERPROOF_SECP160K1_SHA256_SV
`define WYCHERPROOF_SECP160K1_SHA256_SV
typedef struct packed {
  int            tc_id;
  bit            valid;   // Wycheproof: valid/acceptable=1, else=0
  logic [511:0]  hash;    // 固定宣告 512 bits
  logic [527:0]  x;       // 固定宣告 528 bits
  logic [527:0]  y;       // 固定宣告 528 bits
  logic [527:0]  r;       // 固定宣告 528 bits
  logic [527:0]  s;       // 固定宣告 528 bits
} ecdsa_vector_secp160k1_sha256;

localparam int TEST_VECTORS_SECP160K1_SHA256_NUM = 62;

ecdsa_vector_secp160k1_sha256 test_vectors_secp160k1_sha256 [] = '{
  '{2, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'ha89cf5aa14f3e5d8a02f7021c6d0291e7154df23, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{117, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 0, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=0b(0B), s=160b(20B)
  '{125, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h00a89cf5aa14f3e5d8a02f7021c6d0291e7154df, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{133, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=160b(20B)
  '{137, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'ha89cf5aa14f3e5d8a02db727aff07d83a73e2870, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{139, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h57630a55eb0c1a275fd248d8500f827c58c1d790, 160'h1fcb73dfeefa68711c561ca3b9e6056868713540},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{150, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{151, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{152, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h00, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{160, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{161, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{162, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'h01, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{170, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 8'h00},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{171, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 8'h01},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{172, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 8'hff, 8'hff},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{241, 1'b1, 256'h7300000000213f2a525c6035725235c2f696ad3ebb5ee47f140697ad25770d91, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h2e63b73510882b93c69a8d00767f9b9897262b2d, 160'h2e401df2d03607e9a26e16f9550abbc4d40e888c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{242, 1'b1, 256'hddf2000000005e0be0635b245f0b97978afd25daadeb3edb4a0161c27fe06045, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h4296974dca1d2ac6db892b65e2ae5877ab243e1f, 160'h35b0559258b7be92dfa2575d78c9798058e16a4e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{244, 1'b1, 256'ha2bf09460000000076d7dbeffe125eaf02095dff252ee905e296b6350fc311cf, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h0766ca1cad1e6e47a3dc8d86d8ccc18624498273, 160'h47791918c5bb5511cf25194fd52d7cca97a931b5},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{245, 1'b1, 256'h3554e827c700000000e1e75e624a06b3a0a353171160858129e15c544e4f0e65, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h71637fa756fcbc3b8313501c1e651569733ee71a, 160'h12334122b218782a145446996546bcca95c7c968},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{250, 1'b1, 256'h660570d323e9f75fa734000000008792d65ce93eabb7d60d8d9c1bbdcb5ef305, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h6cbe031b8dfd5142eb7c8f69c9d4d3f25f48a903, 160'h27685c54fd837ac971f198b661620eac851d9d7a},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{256, 1'b1, 256'h9ea6994f1e0384c8599aa02e6cf66d9c000000004d89ef50b7e9eb0cfbff7363, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h5b58249bb9fc858db67257a4bb5d21df6d8a1dc5, 160'h74d16dbf41fd4d5bd148a0cc020f6ea6bed1d5eb},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{257, 1'b1, 256'hd03215a8401bcf16693979371a01068a4700000000e2fa5bf692bc670905b18c, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h46fa4b37d994ede647aa00e8552867a0fd932c25, 160'h75a0850d1e7d0d0e3a796a1df069d5bb9eec7309},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{264, 1'b1, 256'he02716d01fb23a5a0068399bf01bab42ef17c6d96e13846c00000000afc0f89d, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h30894ccb595c048cb6ff9dcc5b974b5a72e9fb95, 160'h1c3b805772e98845dbc660d3675174e9842c7f2b},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{265, 1'b1, 256'h9eb0bf583a1a6b9a194e9a16bc7dab2a9061768af89d00659a00000000fc7de1, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h6de326ca60d74a5997d4137b4b6f66f9a6ebff91, 160'h6a5f5b88569920c4f7644a476280a6e711ddf058},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{272, 1'b1, 256'h641227ffffffff6f1b96fa5f097fcf3cc1a3c256870d45a67b83d0967d4b20c0, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h39f9b38cd943bcc3ca0d47a276c419e1ae94643e, 160'h59027aff40966014bdf62c7f6ff1197e5093644c},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{284, 1'b1, 256'h422e82a3d56ed10a9cc21d31d37a25ffffffff67edf7c40204caae73ab0bc75a, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h1c77e9430c235c33a93d7f74ae2b1b67afb75191, 160'h4b1b6c4c49ad002a1017e5017fc495a4ecc85c1e},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{285, 1'b1, 256'h7075d245ccc3281b6e7b329ff738fbb417a5ffffffffa0842d9890b5cf95d018, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h2d3a0bba220b15814b0cac3f1a344f648755ff8e, 160'h68f067f05edd4b543a0d8a92f5a6025769617029},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{287, 1'b1, 256'hde21754e29b85601980bef3d697ea2770ce891a8cdffffffffc7906aa794b39b, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h3174c392114a6e623a4778bbd26dcb8ffd0a5e06, 160'h3425b221031c23d6a99efa813109e53fe5402176},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{290, 1'b1, 256'hfc28259702a03845b6d75219444e8b43d094586e249c8699ffffffffe852512e, 168'h00be74d8dd1d5654265384f74227ab0f8534b5a4fe, 160'h2ab8e5bfeff929794d8dd9c2e3be40e6cf49ad49, 160'h16771ee4085694c00ee10b616484d87e878554d8, 160'h67dffce5c711eca8e370d2bdce36aa0205e7d313},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{299, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h012a78f3ceb2c5606f824b90b4151a7cd788c3c8, 160'h6216521c8b038e7080bb5601ac8b49e96826368b, 8'h03, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=8b(1B), s=8b(1B)
  '{300, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00cee7f5abdb03bb603a30a7a781d2249708931e28, 168'h00f459dfe37fef1cc13d5832452381cc179e708728, 8'h03, 8'h03},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{301, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h48c7400e22d2ef7354b820eb662105e1b6e44a60, 168'h00a329f8bd69afd5aa91d4e18d3cfa2428930dee68, 8'h03, 8'h04},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=8b(1B), s=8b(1B)
  '{305, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h079fdc2ba58d2ce63611b3459035261405e179db, 168'h00dc027bf8924259b02fc4aa144b7dcb58e60eb365, 56'h2d9b4d347952cc, 160'h415936395bb46f9943914f2100607aec6cf33d9d},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=56b(7B), s=160b(20B)
  '{306, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00990cfd22fb6aacfd6cf03761c7e57aa2a5d777d8, 160'h5fce9841ca3a588d3a475e079971814d3ae9fa44, 104'h1033e67e37b32b445580bf4efb, 160'h6b946b946b946b946b9524e49d0953123b068e85},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=104b(13B), s=160b(20B)
  '{310, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6b54692483b37d1cb63c0ba6b5c74af4fbb5b336, 160'h67ea2957b75513d2ae6d1a2ea9ece586da947c9b, 160'h55555555555555555555e8535cf5393398b23ce7, 8'h01},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{311, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h6b54692483b37d1cb63c0ba6b5c74af4fbb5b336, 160'h67ea2957b75513d2ae6d1a2ea9ece586da947c9b, 160'h55555555555555555555e8535cf5393398b23ce7, 8'h00},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=8b(1B)
  '{317, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h41f3d434600a3f8a8a31aebe2cddfe2bc2b0d6e3, 160'h133cd88bbc0a4d81603015f3dce1ea82e1fa49dd, 160'h55555555555555555555e8535cf5393398b23ce3, 160'h55555555555555555555e8535cf5393398b23ce3},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{319, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c1ba77b68c24397599f5eebc6b4a48f4f8caf4c5, 160'h3786ae759de63750382753b333576f5c1b26c540, 40'h0100005383, 160'h7ce6e1f81fbdb6ebf382414e62c1c14200249a82},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{320, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h28a2173e9bcd94c46d5dd3d160c8d3c6f5f392cb, 160'h77ebe984b44814ef24d6d2570ecbea704bf587a0, 40'h0100005383, 160'h2e5c5c1b387dfb0e98740c28008998e351483cfe},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{321, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00fb75a1a2c846d22d787e73d1d7bc7c81b27ce6d4, 160'h4f5ca24aeedd2e6dc1ed2c55f59ef00ce44f800e, 40'h0100005383, 160'h34a4abe436ec3fc4d118f7aceec0df6fdae800d0},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{323, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b5594d926de21168b0f60962e720c7623563158e, 160'h47a500835967a864bcd75d14ae3780ca0f154895, 40'h0100005383, 160'h36155015c2560894b5a1d735e4fe734ef48690c7},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{324, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2df812587ffa67e82da47bce7b72446b7235ea74, 168'h009569210bcbb40d4fd9ce06d58f74b8ecc964bdfb, 40'h0100005383, 160'h6c2aa02b84ac11296b43ae6bc9fce69de90d218e},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{325, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00e3011e8fb90bfdf17424d59d0f7c9757e0a9ba8c, 168'h00ab28c585258001594b87d83dea00294c4a4ee79e, 40'h0100005383, 160'h015c2560894b5a17a0c6dd93d9d5492d33928391},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{326, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c2fb0180784a8f5074304cb708002635e844b3d5, 168'h00c8eff920e00d4ba506c58ca250fcf641b18e6f61, 40'h0100005383, 160'h18f90d4fad917e9601713c4ea95ad2def7b0806f},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{329, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h3943713524548260c840a4c833091e2682bac598, 160'h05acb1d6bca1c685ed1bca4d05dc6ecfb8f22206, 40'h0100005383, 160'h44a5ad0bd0636d9e12be570482bd09b7c9dfcef0},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{330, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h4c21a2c434cac9188f48721e1d0b160d5e3d8502, 160'h73d7e1ccd671a4f7ad0b9b150d4c64a2982191a6, 40'h0100005383, 160'h1a5255f21b761fe2688c7bd677606fb7ed740068},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{331, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h2d36e6f01f0646f272289d73500e4a2fb7450294, 160'h5500bc561c648880fe99476b80b19cc3dfa3169f, 40'h0100005383, 160'h55555555555555555555e8535cf53933ee07ae12},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{332, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h633842757a9dc3b198de959bc34cc10ac9539be2, 160'h14b55c72f731cbec1a6cc80c30c9a868dee85233, 40'h0100005383, 160'h49714251df3ec8f3a9f5a39c44e3be5e5fbfdec4},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{333, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h03688c836288d11d9978ac2cd41ed4884e074555, 160'h1d524a23c8b8871191dee13b6ed4b3dc8ba20105, 40'h0100005383, 160'h599e266b8075ef551833f964e68b1787c9a5d565},  // lens: hash=256b(32B), x=160b(20B), y=160b(20B), r=40b(5B), s=160b(20B)
  '{334, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h37bafb3cba163d05559ca3639906d764b3a213ba, 168'h00b30c713077a32dec18465e1e73568066bef58532, 40'h0100005383, 160'h77f11661e51ad7f10000ce9b8a9fa0b557fdb532},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{335, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c66d00b9cd6b5b5903b2ece209470e712b96f515, 168'h00c9748522a17b59a60e74c69d7de161a5f9ffb532, 40'h0100005383, 160'h11661e51ad7f100000001df88363f82efb0f9833},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{336, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00fe4479b039c9781af875e51a40a1988f99e4777b, 168'h00d4b01aa8430b9a6b271ed609cbe59ad97f189bf5, 40'h0100005383, 160'h22cc3ca35afe200000003bf106c7f05df61f3066},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=40b(5B), s=160b(20B)
  '{345, 1'b0, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h0098defbbf1a0a86d2cfee186065c697f65f471f99, 168'h00e186edcd9ae13a68a8f3030691b2ab20a8b418c6, 160'h55555555555555555555e8535cf5393398b23ce6, 160'h333333333333333333338b6537c655855b9e248a},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{346, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00d3cf5669d7a6aa345133a0ff9f56a88c995a340d, 168'h0094f884562ce27b0b67e0e80e486c4d4e2264e651, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h55555555555555555555e8535cf5393398b23ce6},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{347, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c2e0b6b5d370f374f3b2f5a2e4a01e2bf3c2e158, 160'h5f6879f63a40a9cacc8343214ec2925c47f1d18a, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h49249249249249249249a29098d23107a7743433},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{348, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00b43dd1c55ca1a5af0e9ef4f3b3d30c70feca6f4d, 160'h4fdc2b3171e117fc3e058b7d0ba8818f977ca6d4, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h333333333333333333338b6537c655855b9e248a},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{351, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00862e2eb41fa97389e6d9a5809f33c476255e851c, 160'h6c97ca144a98c842e706d73431d90a366dfcac6a, 160'h74fc71cb95e965fc54ee5fa0227aff946533a0e3, 160'h0eb020c9b97c56649802d1e8ce928dc660acbae8},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{352, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a896b2ce7de0dc53d813053a64a45053f9e6341c, 168'h008f3b7c374dc223c0ff5e32cfc517856ae25ada3e, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h55555555555555555555e8535cf5393398b23ce6},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{353, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00a6b2f424d53ab1dce8ded84894b7c935daa2d869, 160'h576c5baac08c1c5ff45e2b4f5e2c743e24661c7d, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h49249249249249249249a29098d23107a7743433},  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
  '{354, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 160'h299d0559bcd39fb4a5287989d5a02a93ea21db17, 168'h00dc64a6f176f66233d1ccb92bcdde100d39793cd4, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h333333333333333333338b6537c655855b9e248a},  // lens: hash=256b(32B), x=160b(20B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{357, 1'b1, 256'hbb5a52f42f9c9261ed4361f59422a1e30036e7c32b270c8807a419feca605023, 168'h00c05720b3bd92b0f8c72bf85c0772166217234020, 168'h0083a1a12194eda0a5aa53f17f7bff65d6bf5fbb08, 160'h3b4c382ce37aa192a4019e763036f4f5dd4d7ebb, 160'h0eb020c9b97c56649802d1e8ce928dc660acbae8},  // lens: hash=256b(32B), x=168b(21B), y=168b(21B), r=160b(20B), s=160b(20B)
  '{362, 1'b1, 256'he3b0c44298fc1c149afbf4c8996fb92427ae41e4649b934ca495991b7852b855, 168'h008c8b7f800bc9c5588b4970e7559eca926fa38e7b, 160'h6c5d8223426e1cf8d2a2791ab710a14305048ad3, 160'h2e3567b523f24421cf59dc80925775b148eb5380, 160'h38aa38f17c131f0128af4dcafe01e68305414586}  // lens: hash=256b(32B), x=168b(21B), y=160b(20B), r=160b(20B), s=160b(20B)
};
`endif // WYCHERPROOF_SECP160K1_SHA256_SV
